-- Version: v11.9 SP2 11.9.2.1
-- File used only for Simulation

library ieee;
use ieee.std_logic_1164.all;
library smartfusion;
use smartfusion.all;

entity Top is

    port( MSS_RESET_N : in    std_logic;
          SPI_0_DI    : in    std_logic;
          UART_0_RXD  : in    std_logic;
          RD          : out   std_logic_vector(7 downto 0);
          SPI_0_DO    : out   std_logic;
          UART_0_TXD  : out   std_logic;
          SPI_0_CLK   : inout std_logic := 'Z';
          SPI_0_SS    : inout std_logic := 'Z'
        );

end Top;

architecture DEF_ARCH of Top is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DLN1
    port( D : in    std_logic := 'U';
          G : in    std_logic := 'U';
          Q : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOTRI_OB_EB
    port( D    : in    std_logic := 'U';
          E    : in    std_logic := 'U';
          DOUT : out   std_logic;
          EOUT : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AX1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MSS_IF
    port( PIN4    : in    std_logic := 'U';
          PIN5    : in    std_logic := 'U';
          PIN6    : in    std_logic := 'U';
          PIN1    : out   std_logic;
          PIN2    : out   std_logic;
          PIN3    : out   std_logic;
          PIN4INT : out   std_logic;
          PIN5INT : out   std_logic;
          PIN6INT : out   std_logic;
          PIN1INT : in    std_logic := 'U';
          PIN2INT : in    std_logic := 'U';
          PIN3INT : in    std_logic := 'U'
        );
  end component;

  component BUFF
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MSS_APB_IP
    generic (ACT_CONFIG:integer := 0; ACT_FCLK:integer := 0; 
        ACT_DIE:string := ""; ACT_PKG:string := "");

    port( FCLK           : in    std_logic := 'U';
          MACCLKCCC      : in    std_logic := 'U';
          RCOSC          : in    std_logic := 'U';
          MACCLK         : in    std_logic := 'U';
          PLLLOCK        : in    std_logic := 'U';
          MSSRESETn      : in    std_logic := 'U';
          GPOE           : out   std_logic_vector(31 downto 0);
          SPI0DO         : out   std_logic;
          SPI0DOE        : out   std_logic;
          SPI0DI         : in    std_logic := 'U';
          SPI0CLKI       : in    std_logic := 'U';
          SPI0CLKO       : out   std_logic;
          SPI0MODE       : out   std_logic;
          SPI0SSI        : in    std_logic := 'U';
          SPI0SSO        : out   std_logic_vector(7 downto 0);
          UART0TXD       : out   std_logic;
          UART0RXD       : in    std_logic := 'U';
          I2C0SDAI       : in    std_logic := 'U';
          I2C0SDAO       : out   std_logic;
          I2C0SCLI       : in    std_logic := 'U';
          I2C0SCLO       : out   std_logic;
          SPI1DO         : out   std_logic;
          SPI1DOE        : out   std_logic;
          SPI1DI         : in    std_logic := 'U';
          SPI1CLKI       : in    std_logic := 'U';
          SPI1CLKO       : out   std_logic;
          SPI1MODE       : out   std_logic;
          SPI1SSI        : in    std_logic := 'U';
          SPI1SSO        : out   std_logic_vector(7 downto 0);
          UART1TXD       : out   std_logic;
          UART1RXD       : in    std_logic := 'U';
          I2C1SDAI       : in    std_logic := 'U';
          I2C1SDAO       : out   std_logic;
          I2C1SCLI       : in    std_logic := 'U';
          I2C1SCLO       : out   std_logic;
          MACTXD         : out   std_logic_vector(1 downto 0);
          MACRXD         : in    std_logic_vector(1 downto 0) := (others => 'U');
          MACTXEN        : out   std_logic;
          MACCRSDV       : in    std_logic := 'U';
          MACRXER        : in    std_logic := 'U';
          MACMDI         : in    std_logic := 'U';
          MACMDO         : out   std_logic;
          MACMDEN        : out   std_logic;
          MACMDC         : out   std_logic;
          EMCCLK         : out   std_logic;
          EMCCLKRTN      : in    std_logic := 'U';
          EMCRDB         : in    std_logic_vector(15 downto 0) := (others => 'U');
          EMCAB          : out   std_logic_vector(25 downto 0);
          EMCWDB         : out   std_logic_vector(15 downto 0);
          EMCRWn         : out   std_logic;
          EMCCS0n        : out   std_logic;
          EMCCS1n        : out   std_logic;
          EMCOEN0n       : out   std_logic;
          EMCOEN1n       : out   std_logic;
          EMCBYTEN       : out   std_logic_vector(1 downto 0);
          EMCDBOE        : out   std_logic;
          ADC0           : in    std_logic := 'U';
          ADC1           : in    std_logic := 'U';
          ADC2           : in    std_logic := 'U';
          ADC3           : in    std_logic := 'U';
          ADC4           : in    std_logic := 'U';
          ADC5           : in    std_logic := 'U';
          ADC6           : in    std_logic := 'U';
          ADC7           : in    std_logic := 'U';
          ADC8           : in    std_logic := 'U';
          ADC9           : in    std_logic := 'U';
          ADC10          : in    std_logic := 'U';
          ADC11          : in    std_logic := 'U';
          SDD0           : out   std_logic;
          SDD1           : out   std_logic;
          SDD2           : out   std_logic;
          ABPS0          : in    std_logic := 'U';
          ABPS1          : in    std_logic := 'U';
          ABPS2          : in    std_logic := 'U';
          ABPS3          : in    std_logic := 'U';
          ABPS4          : in    std_logic := 'U';
          ABPS5          : in    std_logic := 'U';
          ABPS6          : in    std_logic := 'U';
          ABPS7          : in    std_logic := 'U';
          ABPS8          : in    std_logic := 'U';
          ABPS9          : in    std_logic := 'U';
          ABPS10         : in    std_logic := 'U';
          ABPS11         : in    std_logic := 'U';
          TM0            : in    std_logic := 'U';
          TM1            : in    std_logic := 'U';
          TM2            : in    std_logic := 'U';
          TM3            : in    std_logic := 'U';
          TM4            : in    std_logic := 'U';
          TM5            : in    std_logic := 'U';
          CM0            : in    std_logic := 'U';
          CM1            : in    std_logic := 'U';
          CM2            : in    std_logic := 'U';
          CM3            : in    std_logic := 'U';
          CM4            : in    std_logic := 'U';
          CM5            : in    std_logic := 'U';
          GNDTM0         : in    std_logic := 'U';
          GNDTM1         : in    std_logic := 'U';
          GNDTM2         : in    std_logic := 'U';
          VAREF0         : in    std_logic := 'U';
          VAREF1         : in    std_logic := 'U';
          VAREF2         : in    std_logic := 'U';
          VAREFOUT       : out   std_logic;
          GNDVAREF       : in    std_logic := 'U';
          PUn            : in    std_logic := 'U';
          MSSPADDR       : out   std_logic_vector(19 downto 0);
          MSSPWDATA      : out   std_logic_vector(31 downto 0);
          MSSPRDATA      : in    std_logic_vector(31 downto 0) := (others => 'U');
          FABPADDR       : in    std_logic_vector(31 downto 0) := (others => 'U');
          FABPWDATA      : in    std_logic_vector(31 downto 0) := (others => 'U');
          FABPRDATA      : out   std_logic_vector(31 downto 0);
          DMAREADY       : in    std_logic_vector(1 downto 0) := (others => 'U');
          MSSINT         : out   std_logic_vector(7 downto 0);
          GPI            : in    std_logic_vector(31 downto 0) := (others => 'U');
          GPO            : out   std_logic_vector(31 downto 0);
          MACM2FTXD      : out   std_logic_vector(1 downto 0);
          MACF2MRXD      : in    std_logic_vector(1 downto 0) := (others => 'U');
          ACEFLAGS       : out   std_logic_vector(31 downto 0);
          UART0CTSn      : in    std_logic := 'U';
          UART0DSRn      : in    std_logic := 'U';
          UART0RTSn      : out   std_logic;
          UART0DTRn      : out   std_logic;
          UART0RIn       : in    std_logic := 'U';
          UART0DCDn      : in    std_logic := 'U';
          UART1CTSn      : in    std_logic := 'U';
          UART1DSRn      : in    std_logic := 'U';
          UART1RIn       : in    std_logic := 'U';
          UART1DCDn      : in    std_logic := 'U';
          I2C0SMBALERTNO : out   std_logic;
          I2C0BCLK       : in    std_logic := 'U';
          I2C0SMBALERTNI : in    std_logic := 'U';
          I2C0SMBUSNI    : in    std_logic := 'U';
          I2C1SMBALERTNO : out   std_logic;
          I2C1BCLK       : in    std_logic := 'U';
          I2C1SMBALERTNI : in    std_logic := 'U';
          I2C1SMBUSNI    : in    std_logic := 'U';
          UART1RTSn      : out   std_logic;
          UART1DTRn      : out   std_logic;
          TXEV           : out   std_logic;
          RXEV           : in    std_logic := 'U';
          VRON           : in    std_logic := 'U';
          MACM2FTXEN     : out   std_logic;
          MACF2MCRSDV    : in    std_logic := 'U';
          MACM2FMDEN     : out   std_logic;
          MACF2MRXER     : in    std_logic := 'U';
          MACM2FMDO      : out   std_logic;
          MACF2MMDI      : in    std_logic := 'U';
          MACM2FMDC      : out   std_logic;
          I2C0SMBUSNO    : out   std_logic;
          I2C1SMBUSNO    : out   std_logic;
          CALIBOUT       : out   std_logic;
          CALIBIN        : in    std_logic := 'U';
          LVTTL0         : out   std_logic;
          LVTTL1         : out   std_logic;
          LVTTL2         : out   std_logic;
          LVTTL0EN       : in    std_logic := 'U';
          LVTTL1EN       : in    std_logic := 'U';
          LVTTL2EN       : in    std_logic := 'U';
          LVTTL3         : out   std_logic;
          LVTTL4         : out   std_logic;
          LVTTL5         : out   std_logic;
          LVTTL3EN       : in    std_logic := 'U';
          LVTTL4EN       : in    std_logic := 'U';
          LVTTL5EN       : in    std_logic := 'U';
          LVTTL6         : out   std_logic;
          LVTTL7         : out   std_logic;
          LVTTL8         : out   std_logic;
          LVTTL6EN       : in    std_logic := 'U';
          LVTTL7EN       : in    std_logic := 'U';
          LVTTL8EN       : in    std_logic := 'U';
          LVTTL9         : out   std_logic;
          LVTTL10        : out   std_logic;
          LVTTL11        : out   std_logic;
          LVTTL9EN       : in    std_logic := 'U';
          LVTTL10EN      : in    std_logic := 'U';
          LVTTL11EN      : in    std_logic := 'U';
          CMP0           : out   std_logic;
          CMP1           : out   std_logic;
          CMP2           : out   std_logic;
          CMP3           : out   std_logic;
          CMP4           : out   std_logic;
          CMP5           : out   std_logic;
          FABSDD0D       : in    std_logic := 'U';
          FABSDD1D       : in    std_logic := 'U';
          FABSDD2D       : in    std_logic := 'U';
          CMP6           : out   std_logic;
          CMP7           : out   std_logic;
          CMP8           : out   std_logic;
          FABACETRIG     : in    std_logic := 'U';
          CMP9           : out   std_logic;
          FABSDD0CLK     : in    std_logic := 'U';
          FABSDD1CLK     : in    std_logic := 'U';
          FABSDD2CLK     : in    std_logic := 'U';
          VCC15GOOD      : out   std_logic;
          VCC33GOOD      : out   std_logic;
          PUFABn         : out   std_logic;
          MSSPREADY      : in    std_logic := 'U';
          MSSPSLVERR     : in    std_logic := 'U';
          MSSPSEL        : out   std_logic;
          MSSPENABLE     : out   std_logic;
          MSSPWRITE      : out   std_logic;
          FABPSEL        : in    std_logic := 'U';
          FABPENABLE     : in    std_logic := 'U';
          FABPWRITE      : in    std_logic := 'U';
          FABPREADY      : out   std_logic;
          FABPSLVERR     : out   std_logic;
          DEEPSLEEP      : out   std_logic;
          SLEEP          : out   std_logic;
          M2FRESETn      : out   std_logic;
          WDINT          : out   std_logic;
          FABINT         : in    std_logic := 'U';
          F2MRESETn      : in    std_logic := 'U';
          SYNCCLKFDBK    : in    std_logic := 'U';
          CMP10          : out   std_logic;
          CMP11          : out   std_logic
        );
  end component;

  component DFN1E1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component IOPAD_BI
    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic;
          PAD : inout   std_logic
        );
  end component;

  component IOPAD_TRI
    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IOPAD_IN
    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MSS_CCC_IP
    generic (VCOFREQUENCY:real := 0.0);

    port( CLKA      : in    std_logic := 'U';
          EXTFB     : in    std_logic := 'U';
          GLA       : out   std_logic;
          GLAMSS    : out   std_logic;
          LOCK      : out   std_logic;
          LOCKMSS   : out   std_logic;
          CLKB      : in    std_logic := 'U';
          GLB       : out   std_logic;
          YB        : out   std_logic;
          CLKC      : in    std_logic := 'U';
          GLC       : out   std_logic;
          YC        : out   std_logic;
          MACCLK    : out   std_logic;
          SDIN      : in    std_logic := 'U';
          SCLK      : in    std_logic := 'U';
          SSHIFT    : in    std_logic := 'U';
          SUPDATE   : in    std_logic := 'U';
          MODE      : in    std_logic := 'U';
          SDOUT     : out   std_logic;
          PLLEN     : in    std_logic := 'U';
          OADIV     : in    std_logic_vector(4 downto 0) := (others => 'U');
          OADIVHALF : in    std_logic := 'U';
          OADIVRST  : in    std_logic := 'U';
          OAMUX     : in    std_logic_vector(2 downto 0) := (others => 'U');
          BYPASSA   : in    std_logic := 'U';
          DLYGLA    : in    std_logic_vector(4 downto 0) := (others => 'U');
          DLYGLAMSS : in    std_logic_vector(4 downto 0) := (others => 'U');
          DLYGLAFAB : in    std_logic_vector(4 downto 0) := (others => 'U');
          OBDIV     : in    std_logic_vector(4 downto 0) := (others => 'U');
          OBDIVHALF : in    std_logic := 'U';
          OBDIVRST  : in    std_logic := 'U';
          OBMUX     : in    std_logic_vector(2 downto 0) := (others => 'U');
          BYPASSB   : in    std_logic := 'U';
          DLYGLB    : in    std_logic_vector(4 downto 0) := (others => 'U');
          OCDIV     : in    std_logic_vector(4 downto 0) := (others => 'U');
          OCDIVHALF : in    std_logic := 'U';
          OCDIVRST  : in    std_logic := 'U';
          OCMUX     : in    std_logic_vector(2 downto 0) := (others => 'U');
          BYPASSC   : in    std_logic := 'U';
          DLYGLC    : in    std_logic_vector(4 downto 0) := (others => 'U');
          FINDIV    : in    std_logic_vector(6 downto 0) := (others => 'U');
          FBDIV     : in    std_logic_vector(6 downto 0) := (others => 'U');
          FBDLY     : in    std_logic_vector(4 downto 0) := (others => 'U');
          FBSEL     : in    std_logic_vector(1 downto 0) := (others => 'U');
          XDLYSEL   : in    std_logic := 'U';
          VCOSEL    : in    std_logic_vector(2 downto 0) := (others => 'U');
          GLMUXINT  : in    std_logic := 'U';
          GLMUXSEL  : in    std_logic_vector(1 downto 0) := (others => 'U');
          GLMUXCFG  : in    std_logic_vector(1 downto 0) := (others => 'U')
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKSRC
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MSS_CCC_GL_IF
    port( PIN2    : in    std_logic := 'U';
          PIN3    : in    std_logic := 'U';
          PIN4    : in    std_logic := 'U';
          PIN1    : out   std_logic;
          PIN5    : out   std_logic;
          PIN2INT : out   std_logic;
          PIN3INT : out   std_logic;
          PIN4INT : out   std_logic;
          PIN1INT : in    std_logic := 'U';
          PIN5INT : in    std_logic := 'U'
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MSS_CCC_IF
    port( PIN2    : in    std_logic := 'U';
          PIN3    : in    std_logic := 'U';
          PIN4    : in    std_logic := 'U';
          PIN1    : out   std_logic;
          PIN2INT : out   std_logic;
          PIN3INT : out   std_logic;
          PIN4INT : out   std_logic;
          PIN1INT : in    std_logic := 'U'
        );
  end component;

  component RCOSC
    port( CLKOUT : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port(Y : out std_logic); 
  end component;

  component VCC
    port(Y : out std_logic); 
  end component;

    signal \CoreAPB3_0_APBmslave0_PADDR[0]\, 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, 
        \CoreAPB3_0_APBmslave0_PADDR[5]\, 
        \CoreAPB3_0_APBmslave0_PADDR[6]\, 
        \CoreAPB3_0_APBmslave0_PADDR[7]\, 
        \Intro_0_MSS_MASTER_APB_PADDR[8]\, 
        \Intro_0_MSS_MASTER_APB_PADDR[9]\, 
        \Intro_0_MSS_MASTER_APB_PADDR[10]\, 
        \Intro_0_MSS_MASTER_APB_PADDR[11]\, 
        CoreAPB3_0_APBmslave0_PWRITE, 
        CoreAPB3_0_APBmslave0_PENABLE, 
        Intro_0_MSS_MASTER_APB_PSELx, 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[8]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[9]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[10]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[11]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[12]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[13]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[14]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[15]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[16]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[17]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[18]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[19]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[20]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[21]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[22]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[23]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[24]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[25]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[26]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[27]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[28]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[29]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[30]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[31]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[0]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[1]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[2]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[3]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[4]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[5]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[6]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[7]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[8]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[9]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[10]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[11]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[12]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[13]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[14]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[15]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[16]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[17]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[18]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[19]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[20]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[21]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[22]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[23]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[24]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[25]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[26]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[27]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[28]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[29]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[30]\, 
        \Intro_0_MSS_MASTER_APB_PRDATA[31]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[0]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[1]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[2]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[3]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[4]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[5]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[6]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[7]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[8]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[9]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[10]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[11]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[12]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[13]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[14]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[15]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[16]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[17]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[18]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[19]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[20]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[21]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[22]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[23]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[24]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[25]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[26]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[27]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[28]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[29]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[30]\, 
        \CoreAPB3_0_APBmslave1_PRDATA[31]\, FAB_CLK, 
        Intro_0_M2F_RESET_N, \CoreTimer_0.N_10\, 
        \CoreTimer_0.N_258\, \RD_c[0]\, \RD_c[1]\, \RD_c[2]\, 
        \RD_c[3]\, \RD_c[4]\, \RD_c[5]\, \RD_c[6]\, \RD_c[7]\, 
        \CoreAPB3_0.iPSELS_raw_0[1]\, 
        \CoreAPB3_0.iPSELS_raw_1[1]\, 
        \CoreAPB3_0_APBmslave0_PADDR_0[3]\, 
        \CoreAPB3_0_APBmslave0_PADDR_0[2]\, 
        \Intro_0/MSS_ADLIB_INST_M2FRESETn\, 
        \Intro_0/MSS_UART_0_TXD_D\, \Intro_0/MSS_UART_0_RXD_Y\, 
        \Intro_0/MSS_SPI_0_SS_Y\, \Intro_0/SPI0SSO_net_0[0]\, 
        \Intro_0/MSS_SPI_0_SS_E\, \Intro_0/MSS_SPI_0_DO_D\, 
        \Intro_0/MSS_SPI_0_DO_E\, \Intro_0/MSS_SPI_0_DI_Y\, 
        \Intro_0/MSS_SPI_0_CLK_Y\, \Intro_0/MSS_SPI_0_CLK_D\, 
        \Intro_0/MSS_RESET_0_MSS_RESET_N_Y\, 
        \Intro_0/MSS_ADLIB_INST_EMCCLK\, PLLEN_VCC, GLMUXINT_GND, 
        \Intro_0/GLA0\, \Intro_0/MSS_ADLIB_INST_PLLLOCK\, 
        \Intro_0/MSS_CCC_0/N_CLKA_RCOSC\, 
        \CoreTimer_0/un5_loaden_0\, \CoreTimer_0/N_261\, 
        \CoreTimer_0/Counte_0\, \CoreTimer_0/N_248\, 
        \CoreTimer_0/LoadEnReg_net_1\, 
        \CoreTimer_0/CtrlReg_RNIC1I6A[2]_net_1\, 
        \CoreTimer_0/un1_loadenreg\, 
        \CoreTimer_0/LoadEnReg_RNI42U2A_net_1\, 
        \CoreTimer_0/Count_66_0\, \CoreTimer_0/Count[30]_net_1\, 
        \CoreTimer_0/NextCountPulse_0_0_2\, \CoreTimer_0/N_152\, 
        \CoreTimer_0/NextCountPulse_0_0_a3_0\, 
        \CoreTimer_0/NextCountPulse_0_0_1\, \CoreTimer_0/N_148\, 
        \CoreTimer_0/NextCountPulse_0_0_a3_1_0\, 
        \CoreTimer_0/NextCountPulse_0_0_0\, 
        \CoreTimer_0/NextCountPulse_0_0_a3_2_1\, 
        \CoreTimer_0/N_440\, \CoreTimer_0/N_479\, 
        \CoreTimer_0/NextCountPulse_0_0_a3_4_0\, 
        \CoreTimer_0/TimerPre[1]_net_1\, 
        \CoreTimer_0/TimerPre[2]_net_1\, 
        \CoreTimer_0/PreScale[0]_net_1\, 
        \CoreTimer_0/PreScale[1]_net_1\, 
        \CoreTimer_0/PreScale_n6_i_0_0\, 
        \CoreTimer_0/PreScale_i_0[6]\, \CoreTimer_0/N_150\, 
        \CoreTimer_0/TimerPre[0]_net_1\, 
        \CoreTimer_0/PreScale[7]_net_1\, 
        \CoreTimer_0/TimerPre[3]_net_1\, 
        \CoreTimer_0/PreScale_n2_i_0_0\, 
        \CoreTimer_0/PreScale_i_0[2]\, \CoreTimer_0/N_144\, 
        \CoreTimer_0/PreScale_n4_i_0_0\, 
        \CoreTimer_0/PreScale_i_0[4]\, \CoreTimer_0/N_146\, 
        \CoreTimer_0/PreScale_n3_i_0_0\, 
        \CoreTimer_0/PreScale[3]_net_1\, \CoreTimer_0/N_145\, 
        \CoreTimer_0/PreScale_n5_i_0_0\, 
        \CoreTimer_0/PreScale[5]_net_1\, 
        \CoreTimer_0/PreScale_n8_i_0_a3_0_0_net_1\, 
        \CoreTimer_0/un6_ctrlen_0_a2_0_a2_net_1\, 
        \CoreTimer_0/N_480_1\, \CoreTimer_0/Countlde_0_0_a3_0\, 
        \CoreTimer_0/CountPulse_net_1\, 
        \CoreTimer_0/CtrlReg[0]_net_1\, 
        \CoreTimer_0/N_58_i_0_o2_27\, 
        \CoreTimer_0/N_58_i_0_o2_20\, 
        \CoreTimer_0/N_58_i_0_o2_19\, 
        \CoreTimer_0/N_58_i_0_o2_25\, 
        \CoreTimer_0/N_58_i_0_o2_14\, 
        \CoreTimer_0/N_58_i_0_o2_13\, \CoreTimer_0/N_154\, 
        \CoreTimer_0/N_58_i_0_o2_23\, \CoreTimer_0/N_58_i_0_o2_6\, 
        \CoreTimer_0/N_58_i_0_o2_5\, \CoreTimer_0/N_58_i_0_o2_18\, 
        \CoreTimer_0/N_58_i_0_o2_22\, \CoreTimer_0/N_58_i_0_o2_2\, 
        \CoreTimer_0/N_58_i_0_o2_1\, \CoreTimer_0/N_58_i_0_o2_16\, 
        \CoreTimer_0/Count[28]_net_1\, 
        \CoreTimer_0/Count[29]_net_1\, 
        \CoreTimer_0/N_58_i_0_o2_12\, 
        \CoreTimer_0/Count[21]_net_1\, 
        \CoreTimer_0/Count[18]_net_1\, 
        \CoreTimer_0/N_58_i_0_o2_10\, 
        \CoreTimer_0/Count[23]_net_1\, 
        \CoreTimer_0/Count[9]_net_1\, \CoreTimer_0/N_58_i_0_o2_8\, 
        \CoreTimer_0/Count[4]_net_1\, 
        \CoreTimer_0/Count[8]_net_1\, \CoreTimer_0/N_58_i_0_o2_4\, 
        \CoreTimer_0/Count[24]_net_1\, 
        \CoreTimer_0/Count[31]_net_1\, 
        \CoreTimer_0/Count[25]_net_1\, 
        \CoreTimer_0/Count[10]_net_1\, 
        \CoreTimer_0/Count[11]_net_1\, 
        \CoreTimer_0/Count[20]_net_1\, 
        \CoreTimer_0/Count[22]_net_1\, 
        \CoreTimer_0/Count[16]_net_1\, 
        \CoreTimer_0/Count[19]_net_1\, 
        \CoreTimer_0/Count[17]_net_1\, 
        \CoreTimer_0/Count[15]_net_1\, 
        \CoreTimer_0/Count[13]_net_1\, 
        \CoreTimer_0/Count[7]_net_1\, 
        \CoreTimer_0/Count[3]_net_1\, 
        \CoreTimer_0/Count[5]_net_1\, 
        \CoreTimer_0/Count[6]_net_1\, 
        \CoreTimer_0/Count[14]_net_1\, 
        \CoreTimer_0/Count[12]_net_1\, 
        \CoreTimer_0/Count[26]_net_1\, 
        \CoreTimer_0/Count[27]_net_1\, 
        \CoreTimer_0/NextCountPulse_0_0_a3_0_0\, 
        \CoreTimer_0/PrdataNext_iv_0_i_4[0]\, \CoreTimer_0/N_487\, 
        \CoreTimer_0/N_492\, \CoreTimer_0/N_485\, 
        \CoreTimer_0/PrdataNext_iv_0_i_3[0]\, 
        \CoreTimer_0/Count[0]_net_1\, 
        \CoreTimer_0/PrdataNext_iv_0_i_a3_3_0[0]\, 
        \CoreTimer_0/PrdataNext_iv_0_i_1[0]\, \CoreTimer_0/N_102\, 
        \CoreTimer_0/N_489\, 
        \CoreTimer_0/PrdataNext_0_iv_0_i_1[3]\, 
        \CoreTimer_0/N_151\, \CoreTimer_0/N_257\, 
        \CoreTimer_0/N_244\, 
        \CoreTimer_0/PrdataNext_0_iv_0_i_1[2]\, 
        \CoreTimer_0/Load[2]_net_1\, \CoreTimer_0/N_237\, 
        \CoreTimer_0/PrdataNext_0_iv_0_i_0[2]\, 
        \CoreTimer_0/CtrlReg[2]_net_1\, 
        \CoreTimer_0/PrdataNext_0_iv_0_i_1[1]\, 
        \CoreTimer_0/CtrlReg[1]_net_1\, 
        \CoreTimer_0/iPRDATA_RNO_3[1]_net_1\, 
        \CoreTimer_0/PrdataNext_0_iv_0_i_0[1]\, 
        \CoreTimer_0/Load[1]_net_1\, 
        \CoreTimer_0/un5_intclren_0_a3_0_a3_1\, 
        \CoreTimer_0/N_25\, \CoreTimer_0/N_486\, 
        \CoreTimer_0/IntClr_RNO_net_1\, \CoreTimer_0/N_448\, 
        \CoreTimer_0/N_180\, \CoreTimer_0/Counte\, 
        \CoreTimer_0/N_136\, \CoreTimer_0/N_441\, 
        \CoreTimer_0/PreScale[9]_net_1\, \CoreTimer_0/N_16_2\, 
        \CoreTimer_0/NextCountPulse\, \CoreTimer_0/N_483\, 
        \CoreTimer_0/N_482\, \CoreTimer_0/N_30\, 
        \CoreTimer_0/N_28\, \CoreTimer_0/N_26\, 
        \CoreTimer_0/N_24\, \CoreTimer_0/N_22\, 
        \CoreTimer_0/N_20\, \CoreTimer_0/N_18\, 
        \CoreTimer_0/N_16\, \CoreTimer_0/N_463\, 
        \CoreTimer_0/N_443\, \CoreTimer_0/N_29\, 
        \CoreTimer_0/iPRDATA_RNO_1[1]_net_1\, 
        \CoreTimer_0/iPRDATA_RNO[2]_net_1\, \CoreTimer_0/N_239\, 
        \CoreTimer_0/N_131\, \CoreTimer_0/N_245\, 
        \CoreTimer_0/N_246\, \CoreTimer_0/RawTimInt_RNO_net_1\, 
        \CoreTimer_0/RawTimInt_net_1\, \CoreTimer_0/N_255\, 
        \CoreTimer_0/IntClr_i_0\, \CoreTimer_0/N_385\, 
        \CoreTimer_0/Count_c17\, \CoreTimer_0/N_210\, 
        \CoreTimer_0/N_384\, \CoreTimer_0/Count_c16\, 
        \CoreTimer_0/N_208\, \CoreTimer_0/N_382\, 
        \CoreTimer_0/Count_c14\, \CoreTimer_0/N_204\, 
        \CoreTimer_0/Load[18]_net_1\, 
        \CoreTimer_0/Load[17]_net_1\, 
        \CoreTimer_0/Load[15]_net_1\, \CoreTimer_0/N_393\, 
        \CoreTimer_0/Count_c25\, \CoreTimer_0/N_226\, 
        \CoreTimer_0/N_392\, \CoreTimer_0/Count_c24\, 
        \CoreTimer_0/N_224\, \CoreTimer_0/Count_c26\, 
        \CoreTimer_0/Load[26]_net_1\, 
        \CoreTimer_0/Load[25]_net_1\, \CoreTimer_0/Count_c23\, 
        \CoreTimer_0/Count_c22\, \CoreTimer_0/Count_c18\, 
        \CoreTimer_0/N_447\, \CoreTimer_0/Load[0]_net_1\, 
        \CoreTimer_0/CountIsZeroReg_i_0\, \CoreTimer_0/N_110\, 
        \CoreTimer_0/N_455\, \CoreTimer_0/N_222\, 
        \CoreTimer_0/Load[24]_net_1\, \CoreTimer_0/N_391\, 
        \CoreTimer_0/N_381\, \CoreTimer_0/Count_c13\, 
        \CoreTimer_0/N_202\, \CoreTimer_0/N_379\, 
        \CoreTimer_0/Count_c11\, \CoreTimer_0/N_198\, 
        \CoreTimer_0/Load[14]_net_1\, 
        \CoreTimer_0/Load[12]_net_1\, \CoreTimer_0/N_396\, 
        \CoreTimer_0/Count_c28\, \CoreTimer_0/N_232\, 
        \CoreTimer_0/N_395\, \CoreTimer_0/Count_c27\, 
        \CoreTimer_0/N_230\, \CoreTimer_0/Count_c29\, 
        \CoreTimer_0/Load[29]_net_1\, 
        \CoreTimer_0/Load[28]_net_1\, 
        \CoreTimer_0/PrdataNext[24]\, 
        \CoreTimer_0/DataOut_0_sqmuxa\, \CoreTimer_0/Count_m[24]\, 
        \CoreTimer_0/DataOut_1_sqmuxa\, \CoreTimer_0/Count_c12\, 
        \CoreTimer_0/Count_c15\, 
        \CoreTimer_0/iPRDATA_RNO[12]_net_1\, \CoreTimer_0/N_452\, 
        \CoreTimer_0/N_100\, \CoreTimer_0/N_453\, 
        \CoreTimer_0/N_121\, \CoreTimer_0/N_460\, 
        \CoreTimer_0/N_123\, \CoreTimer_0/N_461\, 
        \CoreTimer_0/PreScale_i_0[8]\, \CoreTimer_0/N_141\, 
        \CoreTimer_0/N_507_mux\, \CoreTimer_0/Counte_mux\, 
        \CoreTimer_0/Count_RNO_1[0]_net_1\, 
        \CoreTimer_0/iPRDATA_RNO_0[30]_net_1\, 
        \CoreTimer_0/Load[30]_net_1\, 
        \CoreTimer_0/iPRDATA_RNO_0[22]_net_1\, 
        \CoreTimer_0/Load[22]_net_1\, 
        \CoreTimer_0/iPRDATA_RNO_0[21]_net_1\, 
        \CoreTimer_0/Load[21]_net_1\, 
        \CoreTimer_0/iPRDATA_RNO_0[20]_net_1\, 
        \CoreTimer_0/Load[20]_net_1\, 
        \CoreTimer_0/iPRDATA_RNO_0[19]_net_1\, 
        \CoreTimer_0/Load[19]_net_1\, 
        \CoreTimer_0/iPRDATA_RNO_0[16]_net_1\, 
        \CoreTimer_0/Load[16]_net_1\, 
        \CoreTimer_0/iPRDATA_RNO_0[8]_net_1\, 
        \CoreTimer_0/Load[8]_net_1\, \CoreTimer_0/N_191_i\, 
        \CoreTimer_0/N_190_i\, \CoreTimer_0/Count[1]_net_1\, 
        \CoreTimer_0/N_153\, \CoreTimer_0/Count[2]_net_1\, 
        \CoreTimer_0/Count_RNO[3]_net_1\, 
        \CoreTimer_0/Load[3]_net_1\, 
        \CoreTimer_0/Count_RNO[1]_net_1\, \CoreTimer_0/N_125\, 
        \CoreTimer_0/N_119\, \CoreTimer_0/N_117\, 
        \CoreTimer_0/N_115\, \CoreTimer_0/N_113\, 
        \CoreTimer_0/N_105\, \CoreTimer_0/N_37\, 
        \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\, 
        \CoreTimer_0/un5_prescaleen_0_a2_1_a3_net_1\, 
        \CoreTimer_0/N_178\, \CoreTimer_0/N_190\, 
        \CoreTimer_0/N_212\, \CoreTimer_0/Count_RNO[2]_net_1\, 
        \CoreTimer_0/Count_RNO[8]_net_1\, \CoreTimer_0/Count_c7\, 
        \CoreTimer_0/Count_RNO[19]_net_1\, 
        \CoreTimer_0/Count_c10\, \CoreTimer_0/Count_c9\, 
        \CoreTimer_0/Count_c8\, \CoreTimer_0/Count_c6\, 
        \CoreTimer_0/Count_c5\, \CoreTimer_0/Count_c4\, 
        \CoreTimer_0/Count_c3\, \CoreTimer_0/Load_m[4]\, 
        \CoreTimer_0/Load[4]_net_1\, \CoreTimer_0/PrdataNext[4]\, 
        \CoreTimer_0/Load_m[6]\, \CoreTimer_0/Load[6]_net_1\, 
        \CoreTimer_0/PrdataNext[6]\, \CoreTimer_0/Load_m[7]\, 
        \CoreTimer_0/Load[7]_net_1\, \CoreTimer_0/PrdataNext[7]\, 
        \CoreTimer_0/N_186\, \CoreTimer_0/N_188\, 
        \CoreTimer_0/Count_RNO[6]_net_1\, 
        \CoreTimer_0/Count_RNO[7]_net_1\, \CoreTimer_0/Load_m[5]\, 
        \CoreTimer_0/Load[5]_net_1\, \CoreTimer_0/PrdataNext[5]\, 
        \CoreTimer_0/Load_m[23]\, \CoreTimer_0/Load[23]_net_1\, 
        \CoreTimer_0/PrdataNext[23]\, \CoreTimer_0/Load_m[25]\, 
        \CoreTimer_0/PrdataNext[25]\, \CoreTimer_0/Load_m[26]\, 
        \CoreTimer_0/PrdataNext[26]\, \CoreTimer_0/Load_m[31]\, 
        \CoreTimer_0/Load[31]_net_1\, 
        \CoreTimer_0/PrdataNext[31]\, \CoreTimer_0/N_182\, 
        \CoreTimer_0/N_184\, \CoreTimer_0/N_192\, 
        \CoreTimer_0/Load[9]_net_1\, \CoreTimer_0/N_194\, 
        \CoreTimer_0/Load[10]_net_1\, \CoreTimer_0/Count_c19\, 
        \CoreTimer_0/N_214\, \CoreTimer_0/Count_c20\, 
        \CoreTimer_0/N_216\, \CoreTimer_0/Count_c21\, 
        \CoreTimer_0/N_218\, \CoreTimer_0/N_220\, 
        \CoreTimer_0/N_228\, \CoreTimer_0/Load[27]_net_1\, 
        \CoreTimer_0/N_234\, \CoreTimer_0/N_236\, 
        \CoreTimer_0/Count_RNO[4]_net_1\, 
        \CoreTimer_0/Count_RNO[5]_net_1\, 
        \CoreTimer_0/Count_RNO[9]_net_1\, 
        \CoreTimer_0/Count_RNO[10]_net_1\, 
        \CoreTimer_0/Count_RNO[20]_net_1\, 
        \CoreTimer_0/Count_RNO[21]_net_1\, 
        \CoreTimer_0/Count_RNO[22]_net_1\, 
        \CoreTimer_0/Count_RNO[23]_net_1\, 
        \CoreTimer_0/Count_RNO[27]_net_1\, 
        \CoreTimer_0/Count_RNO[30]_net_1\, 
        \CoreTimer_0/Count_RNO[31]_net_1\, 
        \CoreTimer_0/Load_m[9]\, \CoreTimer_0/PrdataNext[9]\, 
        \CoreTimer_0/Load_m[10]\, \CoreTimer_0/PrdataNext[10]\, 
        \CoreTimer_0/Load_m[11]\, \CoreTimer_0/Load[11]_net_1\, 
        \CoreTimer_0/PrdataNext[11]\, \CoreTimer_0/Load_m[13]\, 
        \CoreTimer_0/Load[13]_net_1\, 
        \CoreTimer_0/PrdataNext[13]\, \CoreTimer_0/Load_m[15]\, 
        \CoreTimer_0/PrdataNext[15]\, \CoreTimer_0/Load_m[17]\, 
        \CoreTimer_0/PrdataNext[17]\, \CoreTimer_0/Load_m[27]\, 
        \CoreTimer_0/PrdataNext[27]\, \CoreTimer_0/N_196\, 
        \CoreTimer_0/N_200\, \CoreTimer_0/N_206\, 
        \CoreTimer_0/Count_RNO[11]_net_1\, 
        \CoreTimer_0/Count_RNO[13]_net_1\, 
        \CoreTimer_0/Count_RNO[16]_net_1\, 
        \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, 
        \FlashLED_control_wrapper_0/M1/un2_wen_3\, 
        \FlashLED_control_wrapper_0/M1/un2_wen_0\, 
        \FlashLED_control_wrapper_0/M1/un2_wen_1\, 
        \FlashLED_control_wrapper_0/M1/un5_wen_3\, 
        \FlashLED_control_wrapper_0/M1/un5_wen_2\, 
        \FlashLED_control_wrapper_0/M1/un5_wen_1\, 
        \FlashLED_control_wrapper_0/M1/un2_rwclk_5\, 
        \FlashLED_control_wrapper_0/M1/un2_rwclk_3\, 
        \FlashLED_control_wrapper_0/M1/REG_control[5]_net_1\, 
        \FlashLED_control_wrapper_0/M1/REG_control[4]_net_1\, 
        \FlashLED_control_wrapper_0/M1/un2_rwclk_4\, 
        \FlashLED_control_wrapper_0/M1/REG_control[0]_net_1\, 
        \FlashLED_control_wrapper_0/M1/un2_rwclk_1\, 
        \FlashLED_control_wrapper_0/M1/REG_control[1]_net_1\, 
        \FlashLED_control_wrapper_0/M1/REG_control[6]_net_1\, 
        \FlashLED_control_wrapper_0/M1/REG_control[7]_net_1\, 
        \FlashLED_control_wrapper_0/M1/REG_control[2]_net_1\, 
        \FlashLED_control_wrapper_0/M1/REG_control[3]_net_1\, 
        \FlashLED_control_wrapper_0/M1/un2_rwclk\, 
        \FlashLED_control_wrapper_0/M1/un5_wen\, 
        \FlashLED_control_wrapper_0/M1/REG_control_0_sqmuxa_net_1\, 
        \FlashLED_control_wrapper_0/M1/REG_control_1_sqmuxa_net_1\, 
        \FlashLED_control_wrapper_0/M1/REG_load_value[0]_net_1\, 
        \FlashLED_control_wrapper_0/M1/REG_load_value[1]_net_1\, 
        \FlashLED_control_wrapper_0/M1/REG_load_value[2]_net_1\, 
        \FlashLED_control_wrapper_0/M1/REG_load_value[3]_net_1\, 
        \FlashLED_control_wrapper_0/M1/REG_load_value[4]_net_1\, 
        \FlashLED_control_wrapper_0/M1/REG_load_value[5]_net_1\, 
        \FlashLED_control_wrapper_0/M1/REG_load_value[6]_net_1\, 
        \FlashLED_control_wrapper_0/M1/REG_load_value[7]_net_1\, 
        \RD_pad[7]/U0/NET1\, \RD_pad[7]/U0/NET2\, 
        \RD_pad[4]/U0/NET1\, \RD_pad[4]/U0/NET2\, 
        \Intro_0/MSS_CCC_0/I_MSSCCC/SDIN_INT\, 
        \Intro_0/MSS_CCC_0/I_MSSCCC/SCLK_INT\, 
        \Intro_0/MSS_CCC_0/I_MSSCCC/SSHIFT_INT\, 
        \Intro_0/MSS_CCC_0/I_MSSCCC/SDOUT_INT\, 
        \Intro_0/MSS_CCC_0/I_MSSCCC/EXTFB_INT\, 
        \Intro_0/MSS_CCC_0/I_MSSCCC/GLA_INT\, 
        \Intro_0/MSS_CCC_0/I_MSSCCC/LOCK_INT\, 
        \Intro_0/MSS_CCC_0/I_MSSCCC/CLKB_INT\, 
        \Intro_0/MSS_CCC_0/I_MSSCCC/GLB_INT\, 
        \Intro_0/MSS_CCC_0/I_MSSCCC/YB_INT\, 
        \Intro_0/MSS_CCC_0/I_MSSCCC/MODE_INT\, 
        \Intro_0/MSS_CCC_0/I_MSSCCC/CLKC_INT\, 
        \Intro_0/MSS_CCC_0/I_MSSCCC/SUPDATE_INT\, 
        \Intro_0/MSS_CCC_0/I_MSSCCC/GLC_INT\, 
        \Intro_0/MSS_CCC_0/I_MSSCCC/YC_INT\, \RD_pad[2]/U0/NET1\, 
        \RD_pad[2]/U0/NET2\, \RD_pad[5]/U0/NET1\, 
        \RD_pad[5]/U0/NET2\, 
        \Intro_0/MSS_ADLIB_INST/GPO[16]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPO[17]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPO[18]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPI[16]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPI[17]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPI[18]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPO[19]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPO[20]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPO[21]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPI[19]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPI[20]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPI[21]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPO[22]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPO[23]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPO[24]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPI[22]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPI[23]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPI[24]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPO[25]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPO[26]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPO[27]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPI[25]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPI[26]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPI[27]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPO[28]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPO[29]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPO[30]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPI[28]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPI[29]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPI[30]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPO[31]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/SPI0SSO[1]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/SPI0SSO[2]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/GPI[31]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/UART0CTSnINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/UART0DSRnINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/SPI0SSO[3]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/UART0RTSnINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/UART0DTRnINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/UART0RInINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/UART0DCDnINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/UART1CTSnINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/SPI1SSO[1]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/SPI1SSO[2]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/SPI1SSO[3]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/UART1DSRnINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/UART1RInINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/UART1DCDnINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/SPI1SSO[4]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/SPI1SSO[5]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/I2C0SMBALERTNOINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/I2C0BCLKINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/I2C0SMBALERTNIINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/I2C0SMBUSNIINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/SPI1SSO[6]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/SPI1SSO[7]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/I2C1SMBALERTNOINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/I2C1BCLKINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/I2C1SMBALERTNIINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/I2C1SMBUSNIINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/UART1RTSnINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/UART1DTRnINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/TXEVINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/RXEVINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/VRONINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/CALIBININT_NET\, 
        \Intro_0/MSS_ADLIB_INST/I2C0SMBUSNOINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/I2C1SMBUSNOINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/CALIBOUTINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[0]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[1]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[2]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[0]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[1]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[2]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[3]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[4]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[5]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[3]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[4]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[5]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[6]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[7]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[8]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[6]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[7]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[8]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[9]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[10]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[11]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[9]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[10]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[11]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[12]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[13]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[14]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[12]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[13]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[14]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[15]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[16]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[17]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[15]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[16]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[17]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[18]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[19]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[0]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPREADYINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPSLVERRINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[0]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[1]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[2]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[3]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[1]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[2]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[3]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[4]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[5]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[6]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[4]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[5]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[6]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[7]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[8]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[9]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[7]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[8]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[9]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[10]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[11]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[12]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[10]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[11]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[12]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[13]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[14]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[15]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[13]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[14]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[15]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPSELINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPENABLEINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWRITEINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPSELINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPENABLEINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWRITEINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPREADYINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPSLVERRINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/DEEPSLEEPINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[18]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[19]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[20]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/SLEEPINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSINT[0]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSINT[1]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[21]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[22]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[23]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSINT[2]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSINT[3]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSINT[4]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[24]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[25]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[26]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSINT[5]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/M2FRESETnINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSINT[6]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[27]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[28]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[29]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[0]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSINT[7]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/WDINTINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[30]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[31]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[0]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[1]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[2]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[3]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[1]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[2]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[3]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[4]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[5]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[6]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[4]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[5]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[6]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[7]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[8]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[9]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[7]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[8]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[9]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[10]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[11]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[12]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[10]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[11]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[12]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[13]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[14]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[15]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[13]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[14]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[15]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[16]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[17]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[18]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[16]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[17]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[18]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[19]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[20]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[21]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[19]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[20]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[21]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[22]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[23]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[24]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[22]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[23]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[24]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[25]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[26]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[27]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[25]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[26]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[27]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[28]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[29]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[30]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[28]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[29]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[30]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[31]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[31]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABINTINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/F2MRESETnINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/DMAREADY[0]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/DMAREADY[1]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[16]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[17]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[18]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[16]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[17]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[18]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[19]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[20]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[21]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[19]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[20]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[21]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[22]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[23]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[24]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[22]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[23]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[24]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[25]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[26]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[27]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[25]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[26]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[27]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[28]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[29]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[30]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[28]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[29]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[30]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[31]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/SYNCCLKFDBKINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[31]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/LVTTL0INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/LVTTL1INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/LVTTL2INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/LVTTL0ENINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/LVTTL1ENINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/LVTTL2ENINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/LVTTL3INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/LVTTL4INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/LVTTL5INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/LVTTL3ENINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/LVTTL4ENINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/LVTTL5ENINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/LVTTL6INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/LVTTL7INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/LVTTL6ENINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/LVTTL7ENINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/CMP0INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/CMP1INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/CMP2INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/CMP3INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/CMP4INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/CMP5INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABSDD0DINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABSDD1DINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/CMP6INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/CMP7INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABACETRIGINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABSDD0CLKINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/FABSDD1CLKINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[0]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[1]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[2]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[3]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[4]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[5]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[6]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[7]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[8]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[9]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[10]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[11]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[12]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[13]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[14]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[15]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[16]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[17]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[18]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[19]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[20]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[21]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[22]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[23]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[24]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[25]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[26]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[27]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[28]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[29]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[30]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[31]INT_NET\, 
        \Intro_0/MSS_ADLIB_INST/VCC15GOODINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/VCC33GOODINT_NET\, 
        \Intro_0/MSS_ADLIB_INST/PUFABnINT_NET\, 
        \RD_pad[6]/U0/NET1\, \RD_pad[6]/U0/NET2\, 
        \RD_pad[0]/U0/NET1\, \RD_pad[0]/U0/NET2\, 
        \RD_pad[3]/U0/NET1\, \RD_pad[3]/U0/NET2\, 
        \RD_pad[1]/U0/NET1\, \RD_pad[1]/U0/NET2\, AFLSDF_VCC, 
        AFLSDF_GND : std_logic;
    signal GND_power_net1 : std_logic;
    signal VCC_power_net1 : std_logic;
    signal nc47, nc34, nc98, nc89, nc70, nc60, nc74, nc64, nc9, 
        nc92, nc91, nc13, nc23, nc55, nc80, nc33, nc84, nc16, 
        nc26, nc45, nc73, nc58, nc63, nc27, nc17, nc99, nc36, 
        nc48, nc37, nc5, nc101, nc52, nc76, nc51, nc66, nc77, 
        nc67, nc4, nc42, nc100, nc83, nc41, nc90, nc94, nc86, 
        nc59, nc25, nc15, nc87, nc35, nc49, nc28, nc18, nc75, 
        nc65, nc38, nc93, nc1, nc2, nc50, nc22, nc12, nc21, nc11, 
        nc78, nc54, nc68, nc3, nc32, nc40, nc31, nc96, nc44, nc7, 
        nc97, nc85, nc72, nc6, nc71, nc62, nc61, nc19, nc29, nc88, 
        nc53, nc39, nc8, nc82, nc81, nc79, nc43, nc69, nc56, nc20, 
        nc10, nc57, nc95, nc24, nc14, nc46, nc30 : std_logic;

begin 

    GLMUXINT_GND <= GND_power_net1;
    AFLSDF_GND <= GND_power_net1;
    PLLEN_VCC <= VCC_power_net1;
    AFLSDF_VCC <= VCC_power_net1;

    \CoreTimer_0/CountPulse\ : DFN1C0
      port map(D => \CoreTimer_0/NextCountPulse\, CLK => FAB_CLK, 
        CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreTimer_0/CountPulse_net_1\);
    
    \FlashLED_control_wrapper_0/M1/REG_load_value[5]\ : DLN1
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[5]\, G => 
        \FlashLED_control_wrapper_0/M1/REG_control_1_sqmuxa_net_1\, 
        Q => 
        \FlashLED_control_wrapper_0/M1/REG_load_value[5]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO_0[26]\ : NOR2B
      port map(A => \CoreTimer_0/DataOut_0_sqmuxa\, B => 
        \CoreTimer_0/Load[26]_net_1\, Y => 
        \CoreTimer_0/Load_m[26]\);
    
    \CoreTimer_0/iPRDATA_RNO_0[12]\ : MX2
      port map(A => \CoreTimer_0/Load[12]_net_1\, B => 
        \CoreTimer_0/Count[12]_net_1\, S => 
        \CoreAPB3_0_APBmslave0_PADDR_0[2]\, Y => 
        \CoreTimer_0/N_452\);
    
    \RD_pad[3]/U0/U1\ : IOTRI_OB_EB
      port map(D => \RD_c[3]\, E => PLLEN_VCC, DOUT => 
        \RD_pad[3]/U0/NET1\, EOUT => \RD_pad[3]/U0/NET2\);
    
    \CoreTimer_0/PreScale[8]\ : DFN1P0
      port map(D => \CoreTimer_0/N_16\, CLK => FAB_CLK, PRE => 
        Intro_0_M2F_RESET_N, Q => \CoreTimer_0/PreScale_i_0[8]\);
    
    \CoreTimer_0/Load[3]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[3]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0\, Q => 
        \CoreTimer_0/Load[3]_net_1\);
    
    \CoreTimer_0/Count_RNO[28]\ : AX1B
      port map(A => \CoreTimer_0/un1_loadenreg\, B => 
        \CoreTimer_0/Count_c27\, C => \CoreTimer_0/N_230\, Y => 
        \CoreTimer_0/N_395\);
    
    \CoreTimer_0/Count_RNIH5TA5[16]\ : OR2
      port map(A => \CoreTimer_0/Count_c15\, B => 
        \CoreTimer_0/Count[16]_net_1\, Y => 
        \CoreTimer_0/Count_c16\);
    
    \CoreTimer_0/CountPulse_RNO\ : OR3
      port map(A => \CoreTimer_0/N_483\, B => 
        \CoreTimer_0/NextCountPulse_0_0_2\, C => 
        \CoreTimer_0/N_482\, Y => \CoreTimer_0/NextCountPulse\);
    
    \Intro_0/MSS_ADLIB_INST/U_87\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[20]INT_NET\, PIN5INT
         => \Intro_0/MSS_ADLIB_INST/FABPWDATA[19]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/FABPWDATA[21]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[19]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[20]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[21]INT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_47\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[31]INT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[30]INT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[0]INT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[0]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/MSSINT[7]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/WDINTINT_NET\);
    
    \CoreTimer_0/Load[18]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[18]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\, Q => 
        \CoreTimer_0/Load[18]_net_1\);
    
    \CoreTimer_0/Count_RNITBN83[9]\ : OR2
      port map(A => \CoreTimer_0/Count_c8\, B => 
        \CoreTimer_0/Count[9]_net_1\, Y => \CoreTimer_0/Count_c9\);
    
    \Intro_0/MSS_ADLIB_INST_RNIK7F_0\ : BUFF
      port map(A => \CoreAPB3_0_APBmslave0_PADDR[2]\, Y => 
        \CoreAPB3_0_APBmslave0_PADDR_0[2]\);
    
    \CoreTimer_0/Count_RNO[20]\ : AX1B
      port map(A => \CoreTimer_0/Count_c19\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_214\, Y
         => \CoreTimer_0/Count_RNO[20]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO_2[2]\ : AO1A
      port map(A => \CoreTimer_0/Load[2]_net_1\, B => 
        \CoreTimer_0.N_258\, C => \CoreTimer_0/N_237\, Y => 
        \CoreTimer_0/PrdataNext_0_iv_0_i_1[2]\);
    
    \CoreTimer_0/iPRDATA[10]\ : DFN1C0
      port map(D => \CoreTimer_0/PrdataNext[10]\, CLK => FAB_CLK, 
        CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[10]\);
    
    \CoreTimer_0/iPRDATA_RNO_0[25]\ : NOR2B
      port map(A => \CoreTimer_0/DataOut_0_sqmuxa\, B => 
        \CoreTimer_0/Load[25]_net_1\, Y => 
        \CoreTimer_0/Load_m[25]\);
    
    \CoreTimer_0/CountPulse_RNO_5\ : AO1A
      port map(A => \CoreTimer_0/N_148\, B => 
        \CoreTimer_0/NextCountPulse_0_0_a3_1_0\, C => 
        \CoreTimer_0/NextCountPulse_0_0_0\, Y => 
        \CoreTimer_0/NextCountPulse_0_0_1\);
    
    \CoreTimer_0/CtrlReg_RNIC1I6A[2]\ : NOR3B
      port map(A => \CoreTimer_0/CtrlReg[2]_net_1\, B => 
        \CoreTimer_0/PreScale_n8_i_0_a3_0_0_net_1\, C => 
        \CoreTimer_0/N_180\, Y => 
        \CoreTimer_0/CtrlReg_RNIC1I6A[2]_net_1\);
    
    \CoreTimer_0/CtrlReg[0]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[0]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un6_ctrlen_0_a2_0_a2_net_1\, Q => 
        \CoreTimer_0/CtrlReg[0]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO_0[7]\ : NOR2B
      port map(A => \CoreTimer_0/DataOut_0_sqmuxa\, B => 
        \CoreTimer_0/Load[7]_net_1\, Y => \CoreTimer_0/Load_m[7]\);
    
    \Intro_0/MSS_ADLIB_INST/U_58\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => 
        \Intro_0_MSS_MASTER_APB_PRDATA[31]\, PIN6 => GLMUXINT_GND, 
        PIN1 => \CoreAPB3_0_APBmslave0_PWDATA[31]\, PIN2 => OPEN, 
        PIN3 => OPEN, PIN4INT => OPEN, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[31]INT_NET\, PIN6INT
         => OPEN, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[31]INT_NET\, PIN2INT
         => GLMUXINT_GND, PIN3INT => GLMUXINT_GND);
    
    \CoreTimer_0/Count_RNO[11]\ : AX1B
      port map(A => \CoreTimer_0/Count_c10\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_196\, Y
         => \CoreTimer_0/Count_RNO[11]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO_5[0]\ : OR3A
      port map(A => \CoreTimer_0/N_102\, B => 
        CoreAPB3_0_APBmslave0_PWRITE, C => \CoreTimer_0/N_489\, Y
         => \CoreTimer_0/PrdataNext_iv_0_i_1[0]\);
    
    \CoreTimer_0/CountPulse_RNO_11\ : OR2A
      port map(A => \CoreTimer_0/TimerPre[0]_net_1\, B => 
        \CoreTimer_0/PreScale[3]_net_1\, Y => \CoreTimer_0/N_443\);
    
    \CoreTimer_0/CountPulse_RNO_0\ : NOR3A
      port map(A => \CoreTimer_0/NextCountPulse_0_0_a3_4_0\, B
         => \CoreTimer_0/TimerPre[0]_net_1\, C => 
        \CoreTimer_0/N_441\, Y => \CoreTimer_0/N_483\);
    
    \CoreTimer_0/Count_RNO_0[22]\ : MX2
      port map(A => \CoreTimer_0/Count[22]_net_1\, B => 
        \CoreTimer_0/Load[22]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_218\);
    
    \CoreTimer_0/Count_RNIRAUK[5]\ : OR2
      port map(A => \CoreTimer_0/Count[5]_net_1\, B => 
        \CoreTimer_0/Count[6]_net_1\, Y => 
        \CoreTimer_0/N_58_i_0_o2_4\);
    
    \CoreTimer_0/PreScale[0]\ : DFN1C0
      port map(D => \CoreTimer_0/N_141\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => \CoreTimer_0/PreScale[0]_net_1\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_19\ : NOR3C
      port map(A => \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, B => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[19]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[19]\);
    
    \Intro_0/MSS_ADLIB_INST/U_92\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => GLMUXINT_GND, PIN2INT => GLMUXINT_GND, PIN3INT
         => GLMUXINT_GND);
    
    \Intro_0/MSS_ADLIB_INST/U_9\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => \Intro_0/MSS_ADLIB_INST/UART1RInINT_NET\, 
        PIN5INT => \Intro_0/MSS_ADLIB_INST/UART1DSRnINT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/UART1DCDnINT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/SPI1SSO[1]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/SPI1SSO[2]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/SPI1SSO[3]INT_NET\);
    
    \CoreTimer_0/un6_ctrlen_0_a2_0_a2\ : NOR2B
      port map(A => \CoreTimer_0/N_261\, B => \CoreTimer_0/N_257\, 
        Y => \CoreTimer_0/un6_ctrlen_0_a2_0_a2_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_80\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[14]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[15]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[16]INT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_40\ : MSS_IF
      port map(PIN4 => \Intro_0_MSS_MASTER_APB_PRDATA[11]\, PIN5
         => \Intro_0_MSS_MASTER_APB_PRDATA[10]\, PIN6 => 
        \Intro_0_MSS_MASTER_APB_PRDATA[12]\, PIN1 => 
        \CoreAPB3_0_APBmslave0_PWDATA[10]\, PIN2 => 
        \CoreAPB3_0_APBmslave0_PWDATA[11]\, PIN3 => 
        \CoreAPB3_0_APBmslave0_PWDATA[12]\, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[11]INT_NET\, PIN5INT
         => \Intro_0/MSS_ADLIB_INST/MSSPRDATA[10]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/MSSPRDATA[12]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[10]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[11]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[12]INT_NET\);
    
    \FlashLED_control_wrapper_0/M1/REG_control[7]\ : DLN1
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[7]\, G => 
        \FlashLED_control_wrapper_0/M1/REG_control_0_sqmuxa_net_1\, 
        Q => \FlashLED_control_wrapper_0/M1/REG_control[7]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO[24]\ : AO1
      port map(A => \CoreTimer_0/DataOut_0_sqmuxa\, B => 
        \CoreTimer_0/Load[24]_net_1\, C => 
        \CoreTimer_0/Count_m[24]\, Y => 
        \CoreTimer_0/PrdataNext[24]\);
    
    \CoreTimer_0/Count_RNO[17]\ : AX1B
      port map(A => \CoreTimer_0/un1_loadenreg\, B => 
        \CoreTimer_0/Count_c16\, C => \CoreTimer_0/N_208\, Y => 
        \CoreTimer_0/N_384\);
    
    \CoreTimer_0/Count_RNO[16]\ : AX1B
      port map(A => \CoreTimer_0/Count_c15\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_206\, Y
         => \CoreTimer_0/Count_RNO[16]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_CORE\ : MSS_APB_IP
      generic map(ACT_CONFIG => 0, ACT_FCLK => 32000000,
         ACT_DIE => "IP4X3M1", ACT_PKG => "fg484")

      port map(FCLK => \Intro_0/GLA0\, MACCLKCCC => GLMUXINT_GND, 
        RCOSC => GLMUXINT_GND, MACCLK => GLMUXINT_GND, PLLLOCK
         => \Intro_0/MSS_ADLIB_INST_PLLLOCK\, MSSRESETn => 
        \Intro_0/MSS_RESET_0_MSS_RESET_N_Y\, GPOE(31) => nc47, 
        GPOE(30) => nc34, GPOE(29) => nc98, GPOE(28) => nc89, 
        GPOE(27) => nc70, GPOE(26) => nc60, GPOE(25) => nc74, 
        GPOE(24) => nc64, GPOE(23) => nc9, GPOE(22) => nc92, 
        GPOE(21) => nc91, GPOE(20) => nc13, GPOE(19) => nc23, 
        GPOE(18) => nc55, GPOE(17) => nc80, GPOE(16) => nc33, 
        GPOE(15) => nc84, GPOE(14) => nc16, GPOE(13) => nc26, 
        GPOE(12) => nc45, GPOE(11) => nc73, GPOE(10) => nc58, 
        GPOE(9) => nc63, GPOE(8) => nc27, GPOE(7) => nc17, 
        GPOE(6) => nc99, GPOE(5) => nc36, GPOE(4) => nc48, 
        GPOE(3) => nc37, GPOE(2) => nc5, GPOE(1) => nc101, 
        GPOE(0) => nc52, SPI0DO => \Intro_0/MSS_SPI_0_DO_D\, 
        SPI0DOE => \Intro_0/MSS_SPI_0_DO_E\, SPI0DI => 
        \Intro_0/MSS_SPI_0_DI_Y\, SPI0CLKI => 
        \Intro_0/MSS_SPI_0_CLK_Y\, SPI0CLKO => 
        \Intro_0/MSS_SPI_0_CLK_D\, SPI0MODE => 
        \Intro_0/MSS_SPI_0_SS_E\, SPI0SSI => 
        \Intro_0/MSS_SPI_0_SS_Y\, SPI0SSO(7) => nc76, SPI0SSO(6)
         => nc51, SPI0SSO(5) => nc66, SPI0SSO(4) => nc77, 
        SPI0SSO(3) => \Intro_0/MSS_ADLIB_INST/SPI0SSO[3]INT_NET\, 
        SPI0SSO(2) => \Intro_0/MSS_ADLIB_INST/SPI0SSO[2]INT_NET\, 
        SPI0SSO(1) => \Intro_0/MSS_ADLIB_INST/SPI0SSO[1]INT_NET\, 
        SPI0SSO(0) => \Intro_0/SPI0SSO_net_0[0]\, UART0TXD => 
        \Intro_0/MSS_UART_0_TXD_D\, UART0RXD => 
        \Intro_0/MSS_UART_0_RXD_Y\, I2C0SDAI => GLMUXINT_GND, 
        I2C0SDAO => OPEN, I2C0SCLI => GLMUXINT_GND, I2C0SCLO => 
        OPEN, SPI1DO => OPEN, SPI1DOE => OPEN, SPI1DI => 
        GLMUXINT_GND, SPI1CLKI => GLMUXINT_GND, SPI1CLKO => OPEN, 
        SPI1MODE => OPEN, SPI1SSI => GLMUXINT_GND, SPI1SSO(7) => 
        \Intro_0/MSS_ADLIB_INST/SPI1SSO[7]INT_NET\, SPI1SSO(6)
         => \Intro_0/MSS_ADLIB_INST/SPI1SSO[6]INT_NET\, 
        SPI1SSO(5) => \Intro_0/MSS_ADLIB_INST/SPI1SSO[5]INT_NET\, 
        SPI1SSO(4) => \Intro_0/MSS_ADLIB_INST/SPI1SSO[4]INT_NET\, 
        SPI1SSO(3) => \Intro_0/MSS_ADLIB_INST/SPI1SSO[3]INT_NET\, 
        SPI1SSO(2) => \Intro_0/MSS_ADLIB_INST/SPI1SSO[2]INT_NET\, 
        SPI1SSO(1) => \Intro_0/MSS_ADLIB_INST/SPI1SSO[1]INT_NET\, 
        SPI1SSO(0) => nc67, UART1TXD => OPEN, UART1RXD => 
        GLMUXINT_GND, I2C1SDAI => GLMUXINT_GND, I2C1SDAO => OPEN, 
        I2C1SCLI => GLMUXINT_GND, I2C1SCLO => OPEN, MACTXD(1) => 
        nc4, MACTXD(0) => nc42, MACRXD(1) => GLMUXINT_GND, 
        MACRXD(0) => GLMUXINT_GND, MACTXEN => OPEN, MACCRSDV => 
        GLMUXINT_GND, MACRXER => GLMUXINT_GND, MACMDI => 
        GLMUXINT_GND, MACMDO => OPEN, MACMDEN => OPEN, MACMDC => 
        OPEN, EMCCLK => \Intro_0/MSS_ADLIB_INST_EMCCLK\, 
        EMCCLKRTN => \Intro_0/MSS_ADLIB_INST_EMCCLK\, EMCRDB(15)
         => GLMUXINT_GND, EMCRDB(14) => GLMUXINT_GND, EMCRDB(13)
         => GLMUXINT_GND, EMCRDB(12) => GLMUXINT_GND, EMCRDB(11)
         => GLMUXINT_GND, EMCRDB(10) => GLMUXINT_GND, EMCRDB(9)
         => GLMUXINT_GND, EMCRDB(8) => GLMUXINT_GND, EMCRDB(7)
         => GLMUXINT_GND, EMCRDB(6) => GLMUXINT_GND, EMCRDB(5)
         => GLMUXINT_GND, EMCRDB(4) => GLMUXINT_GND, EMCRDB(3)
         => GLMUXINT_GND, EMCRDB(2) => GLMUXINT_GND, EMCRDB(1)
         => GLMUXINT_GND, EMCRDB(0) => GLMUXINT_GND, EMCAB(25)
         => nc100, EMCAB(24) => nc83, EMCAB(23) => nc41, 
        EMCAB(22) => nc90, EMCAB(21) => nc94, EMCAB(20) => nc86, 
        EMCAB(19) => nc59, EMCAB(18) => nc25, EMCAB(17) => nc15, 
        EMCAB(16) => nc87, EMCAB(15) => nc35, EMCAB(14) => nc49, 
        EMCAB(13) => nc28, EMCAB(12) => nc18, EMCAB(11) => nc75, 
        EMCAB(10) => nc65, EMCAB(9) => nc38, EMCAB(8) => nc93, 
        EMCAB(7) => nc1, EMCAB(6) => nc2, EMCAB(5) => nc50, 
        EMCAB(4) => nc22, EMCAB(3) => nc12, EMCAB(2) => nc21, 
        EMCAB(1) => nc11, EMCAB(0) => nc78, EMCWDB(15) => nc54, 
        EMCWDB(14) => nc68, EMCWDB(13) => nc3, EMCWDB(12) => nc32, 
        EMCWDB(11) => nc40, EMCWDB(10) => nc31, EMCWDB(9) => nc96, 
        EMCWDB(8) => nc44, EMCWDB(7) => nc7, EMCWDB(6) => nc97, 
        EMCWDB(5) => nc85, EMCWDB(4) => nc72, EMCWDB(3) => nc6, 
        EMCWDB(2) => nc71, EMCWDB(1) => nc62, EMCWDB(0) => nc61, 
        EMCRWn => OPEN, EMCCS0n => OPEN, EMCCS1n => OPEN, 
        EMCOEN0n => OPEN, EMCOEN1n => OPEN, EMCBYTEN(1) => nc19, 
        EMCBYTEN(0) => nc29, EMCDBOE => OPEN, ADC0 => 
        GLMUXINT_GND, ADC1 => GLMUXINT_GND, ADC2 => GLMUXINT_GND, 
        ADC3 => GLMUXINT_GND, ADC4 => GLMUXINT_GND, ADC5 => 
        GLMUXINT_GND, ADC6 => GLMUXINT_GND, ADC7 => GLMUXINT_GND, 
        ADC8 => GLMUXINT_GND, ADC9 => GLMUXINT_GND, ADC10 => 
        GLMUXINT_GND, ADC11 => GLMUXINT_GND, SDD0 => OPEN, SDD1
         => OPEN, SDD2 => OPEN, ABPS0 => GLMUXINT_GND, ABPS1 => 
        GLMUXINT_GND, ABPS2 => GLMUXINT_GND, ABPS3 => 
        GLMUXINT_GND, ABPS4 => GLMUXINT_GND, ABPS5 => 
        GLMUXINT_GND, ABPS6 => GLMUXINT_GND, ABPS7 => 
        GLMUXINT_GND, ABPS8 => GLMUXINT_GND, ABPS9 => 
        GLMUXINT_GND, ABPS10 => GLMUXINT_GND, ABPS11 => 
        GLMUXINT_GND, TM0 => GLMUXINT_GND, TM1 => GLMUXINT_GND, 
        TM2 => GLMUXINT_GND, TM3 => GLMUXINT_GND, TM4 => 
        GLMUXINT_GND, TM5 => GLMUXINT_GND, CM0 => GLMUXINT_GND, 
        CM1 => GLMUXINT_GND, CM2 => GLMUXINT_GND, CM3 => 
        GLMUXINT_GND, CM4 => GLMUXINT_GND, CM5 => GLMUXINT_GND, 
        GNDTM0 => GLMUXINT_GND, GNDTM1 => GLMUXINT_GND, GNDTM2
         => GLMUXINT_GND, VAREF0 => GLMUXINT_GND, VAREF1 => 
        GLMUXINT_GND, VAREF2 => GLMUXINT_GND, VAREFOUT => OPEN, 
        GNDVAREF => GLMUXINT_GND, PUn => GLMUXINT_GND, 
        MSSPADDR(19) => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[19]INT_NET\, 
        MSSPADDR(18) => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[18]INT_NET\, 
        MSSPADDR(17) => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[17]INT_NET\, 
        MSSPADDR(16) => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[16]INT_NET\, 
        MSSPADDR(15) => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[15]INT_NET\, 
        MSSPADDR(14) => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[14]INT_NET\, 
        MSSPADDR(13) => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[13]INT_NET\, 
        MSSPADDR(12) => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[12]INT_NET\, 
        MSSPADDR(11) => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[11]INT_NET\, 
        MSSPADDR(10) => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[10]INT_NET\, MSSPADDR(9)
         => \Intro_0/MSS_ADLIB_INST/MSSPADDR[9]INT_NET\, 
        MSSPADDR(8) => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[8]INT_NET\, MSSPADDR(7)
         => \Intro_0/MSS_ADLIB_INST/MSSPADDR[7]INT_NET\, 
        MSSPADDR(6) => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[6]INT_NET\, MSSPADDR(5)
         => \Intro_0/MSS_ADLIB_INST/MSSPADDR[5]INT_NET\, 
        MSSPADDR(4) => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[4]INT_NET\, MSSPADDR(3)
         => \Intro_0/MSS_ADLIB_INST/MSSPADDR[3]INT_NET\, 
        MSSPADDR(2) => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[2]INT_NET\, MSSPADDR(1)
         => \Intro_0/MSS_ADLIB_INST/MSSPADDR[1]INT_NET\, 
        MSSPADDR(0) => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[0]INT_NET\, 
        MSSPWDATA(31) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[31]INT_NET\, 
        MSSPWDATA(30) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[30]INT_NET\, 
        MSSPWDATA(29) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[29]INT_NET\, 
        MSSPWDATA(28) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[28]INT_NET\, 
        MSSPWDATA(27) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[27]INT_NET\, 
        MSSPWDATA(26) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[26]INT_NET\, 
        MSSPWDATA(25) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[25]INT_NET\, 
        MSSPWDATA(24) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[24]INT_NET\, 
        MSSPWDATA(23) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[23]INT_NET\, 
        MSSPWDATA(22) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[22]INT_NET\, 
        MSSPWDATA(21) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[21]INT_NET\, 
        MSSPWDATA(20) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[20]INT_NET\, 
        MSSPWDATA(19) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[19]INT_NET\, 
        MSSPWDATA(18) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[18]INT_NET\, 
        MSSPWDATA(17) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[17]INT_NET\, 
        MSSPWDATA(16) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[16]INT_NET\, 
        MSSPWDATA(15) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[15]INT_NET\, 
        MSSPWDATA(14) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[14]INT_NET\, 
        MSSPWDATA(13) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[13]INT_NET\, 
        MSSPWDATA(12) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[12]INT_NET\, 
        MSSPWDATA(11) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[11]INT_NET\, 
        MSSPWDATA(10) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[10]INT_NET\, 
        MSSPWDATA(9) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[9]INT_NET\, 
        MSSPWDATA(8) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[8]INT_NET\, 
        MSSPWDATA(7) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[7]INT_NET\, 
        MSSPWDATA(6) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[6]INT_NET\, 
        MSSPWDATA(5) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[5]INT_NET\, 
        MSSPWDATA(4) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[4]INT_NET\, 
        MSSPWDATA(3) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[3]INT_NET\, 
        MSSPWDATA(2) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[2]INT_NET\, 
        MSSPWDATA(1) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[1]INT_NET\, 
        MSSPWDATA(0) => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[0]INT_NET\, 
        MSSPRDATA(31) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[31]INT_NET\, 
        MSSPRDATA(30) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[30]INT_NET\, 
        MSSPRDATA(29) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[29]INT_NET\, 
        MSSPRDATA(28) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[28]INT_NET\, 
        MSSPRDATA(27) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[27]INT_NET\, 
        MSSPRDATA(26) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[26]INT_NET\, 
        MSSPRDATA(25) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[25]INT_NET\, 
        MSSPRDATA(24) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[24]INT_NET\, 
        MSSPRDATA(23) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[23]INT_NET\, 
        MSSPRDATA(22) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[22]INT_NET\, 
        MSSPRDATA(21) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[21]INT_NET\, 
        MSSPRDATA(20) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[20]INT_NET\, 
        MSSPRDATA(19) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[19]INT_NET\, 
        MSSPRDATA(18) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[18]INT_NET\, 
        MSSPRDATA(17) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[17]INT_NET\, 
        MSSPRDATA(16) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[16]INT_NET\, 
        MSSPRDATA(15) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[15]INT_NET\, 
        MSSPRDATA(14) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[14]INT_NET\, 
        MSSPRDATA(13) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[13]INT_NET\, 
        MSSPRDATA(12) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[12]INT_NET\, 
        MSSPRDATA(11) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[11]INT_NET\, 
        MSSPRDATA(10) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[10]INT_NET\, 
        MSSPRDATA(9) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[9]INT_NET\, 
        MSSPRDATA(8) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[8]INT_NET\, 
        MSSPRDATA(7) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[7]INT_NET\, 
        MSSPRDATA(6) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[6]INT_NET\, 
        MSSPRDATA(5) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[5]INT_NET\, 
        MSSPRDATA(4) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[4]INT_NET\, 
        MSSPRDATA(3) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[3]INT_NET\, 
        MSSPRDATA(2) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[2]INT_NET\, 
        MSSPRDATA(1) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[1]INT_NET\, 
        MSSPRDATA(0) => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[0]INT_NET\, 
        FABPADDR(31) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[31]INT_NET\, 
        FABPADDR(30) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[30]INT_NET\, 
        FABPADDR(29) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[29]INT_NET\, 
        FABPADDR(28) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[28]INT_NET\, 
        FABPADDR(27) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[27]INT_NET\, 
        FABPADDR(26) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[26]INT_NET\, 
        FABPADDR(25) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[25]INT_NET\, 
        FABPADDR(24) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[24]INT_NET\, 
        FABPADDR(23) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[23]INT_NET\, 
        FABPADDR(22) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[22]INT_NET\, 
        FABPADDR(21) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[21]INT_NET\, 
        FABPADDR(20) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[20]INT_NET\, 
        FABPADDR(19) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[19]INT_NET\, 
        FABPADDR(18) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[18]INT_NET\, 
        FABPADDR(17) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[17]INT_NET\, 
        FABPADDR(16) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[16]INT_NET\, 
        FABPADDR(15) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[15]INT_NET\, 
        FABPADDR(14) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[14]INT_NET\, 
        FABPADDR(13) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[13]INT_NET\, 
        FABPADDR(12) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[12]INT_NET\, 
        FABPADDR(11) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[11]INT_NET\, 
        FABPADDR(10) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[10]INT_NET\, FABPADDR(9)
         => \Intro_0/MSS_ADLIB_INST/FABPADDR[9]INT_NET\, 
        FABPADDR(8) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[8]INT_NET\, FABPADDR(7)
         => \Intro_0/MSS_ADLIB_INST/FABPADDR[7]INT_NET\, 
        FABPADDR(6) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[6]INT_NET\, FABPADDR(5)
         => \Intro_0/MSS_ADLIB_INST/FABPADDR[5]INT_NET\, 
        FABPADDR(4) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[4]INT_NET\, FABPADDR(3)
         => \Intro_0/MSS_ADLIB_INST/FABPADDR[3]INT_NET\, 
        FABPADDR(2) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[2]INT_NET\, FABPADDR(1)
         => \Intro_0/MSS_ADLIB_INST/FABPADDR[1]INT_NET\, 
        FABPADDR(0) => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[0]INT_NET\, 
        FABPWDATA(31) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[31]INT_NET\, 
        FABPWDATA(30) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[30]INT_NET\, 
        FABPWDATA(29) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[29]INT_NET\, 
        FABPWDATA(28) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[28]INT_NET\, 
        FABPWDATA(27) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[27]INT_NET\, 
        FABPWDATA(26) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[26]INT_NET\, 
        FABPWDATA(25) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[25]INT_NET\, 
        FABPWDATA(24) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[24]INT_NET\, 
        FABPWDATA(23) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[23]INT_NET\, 
        FABPWDATA(22) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[22]INT_NET\, 
        FABPWDATA(21) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[21]INT_NET\, 
        FABPWDATA(20) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[20]INT_NET\, 
        FABPWDATA(19) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[19]INT_NET\, 
        FABPWDATA(18) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[18]INT_NET\, 
        FABPWDATA(17) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[17]INT_NET\, 
        FABPWDATA(16) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[16]INT_NET\, 
        FABPWDATA(15) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[15]INT_NET\, 
        FABPWDATA(14) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[14]INT_NET\, 
        FABPWDATA(13) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[13]INT_NET\, 
        FABPWDATA(12) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[12]INT_NET\, 
        FABPWDATA(11) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[11]INT_NET\, 
        FABPWDATA(10) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[10]INT_NET\, 
        FABPWDATA(9) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[9]INT_NET\, 
        FABPWDATA(8) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[8]INT_NET\, 
        FABPWDATA(7) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[7]INT_NET\, 
        FABPWDATA(6) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[6]INT_NET\, 
        FABPWDATA(5) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[5]INT_NET\, 
        FABPWDATA(4) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[4]INT_NET\, 
        FABPWDATA(3) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[3]INT_NET\, 
        FABPWDATA(2) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[2]INT_NET\, 
        FABPWDATA(1) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[1]INT_NET\, 
        FABPWDATA(0) => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[0]INT_NET\, 
        FABPRDATA(31) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[31]INT_NET\, 
        FABPRDATA(30) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[30]INT_NET\, 
        FABPRDATA(29) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[29]INT_NET\, 
        FABPRDATA(28) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[28]INT_NET\, 
        FABPRDATA(27) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[27]INT_NET\, 
        FABPRDATA(26) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[26]INT_NET\, 
        FABPRDATA(25) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[25]INT_NET\, 
        FABPRDATA(24) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[24]INT_NET\, 
        FABPRDATA(23) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[23]INT_NET\, 
        FABPRDATA(22) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[22]INT_NET\, 
        FABPRDATA(21) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[21]INT_NET\, 
        FABPRDATA(20) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[20]INT_NET\, 
        FABPRDATA(19) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[19]INT_NET\, 
        FABPRDATA(18) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[18]INT_NET\, 
        FABPRDATA(17) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[17]INT_NET\, 
        FABPRDATA(16) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[16]INT_NET\, 
        FABPRDATA(15) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[15]INT_NET\, 
        FABPRDATA(14) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[14]INT_NET\, 
        FABPRDATA(13) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[13]INT_NET\, 
        FABPRDATA(12) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[12]INT_NET\, 
        FABPRDATA(11) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[11]INT_NET\, 
        FABPRDATA(10) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[10]INT_NET\, 
        FABPRDATA(9) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[9]INT_NET\, 
        FABPRDATA(8) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[8]INT_NET\, 
        FABPRDATA(7) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[7]INT_NET\, 
        FABPRDATA(6) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[6]INT_NET\, 
        FABPRDATA(5) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[5]INT_NET\, 
        FABPRDATA(4) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[4]INT_NET\, 
        FABPRDATA(3) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[3]INT_NET\, 
        FABPRDATA(2) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[2]INT_NET\, 
        FABPRDATA(1) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[1]INT_NET\, 
        FABPRDATA(0) => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[0]INT_NET\, DMAREADY(1)
         => \Intro_0/MSS_ADLIB_INST/DMAREADY[1]INT_NET\, 
        DMAREADY(0) => 
        \Intro_0/MSS_ADLIB_INST/DMAREADY[0]INT_NET\, MSSINT(7)
         => \Intro_0/MSS_ADLIB_INST/MSSINT[7]INT_NET\, MSSINT(6)
         => \Intro_0/MSS_ADLIB_INST/MSSINT[6]INT_NET\, MSSINT(5)
         => \Intro_0/MSS_ADLIB_INST/MSSINT[5]INT_NET\, MSSINT(4)
         => \Intro_0/MSS_ADLIB_INST/MSSINT[4]INT_NET\, MSSINT(3)
         => \Intro_0/MSS_ADLIB_INST/MSSINT[3]INT_NET\, MSSINT(2)
         => \Intro_0/MSS_ADLIB_INST/MSSINT[2]INT_NET\, MSSINT(1)
         => \Intro_0/MSS_ADLIB_INST/MSSINT[1]INT_NET\, MSSINT(0)
         => \Intro_0/MSS_ADLIB_INST/MSSINT[0]INT_NET\, GPI(31)
         => \Intro_0/MSS_ADLIB_INST/GPI[31]INT_NET\, GPI(30) => 
        \Intro_0/MSS_ADLIB_INST/GPI[30]INT_NET\, GPI(29) => 
        \Intro_0/MSS_ADLIB_INST/GPI[29]INT_NET\, GPI(28) => 
        \Intro_0/MSS_ADLIB_INST/GPI[28]INT_NET\, GPI(27) => 
        \Intro_0/MSS_ADLIB_INST/GPI[27]INT_NET\, GPI(26) => 
        \Intro_0/MSS_ADLIB_INST/GPI[26]INT_NET\, GPI(25) => 
        \Intro_0/MSS_ADLIB_INST/GPI[25]INT_NET\, GPI(24) => 
        \Intro_0/MSS_ADLIB_INST/GPI[24]INT_NET\, GPI(23) => 
        \Intro_0/MSS_ADLIB_INST/GPI[23]INT_NET\, GPI(22) => 
        \Intro_0/MSS_ADLIB_INST/GPI[22]INT_NET\, GPI(21) => 
        \Intro_0/MSS_ADLIB_INST/GPI[21]INT_NET\, GPI(20) => 
        \Intro_0/MSS_ADLIB_INST/GPI[20]INT_NET\, GPI(19) => 
        \Intro_0/MSS_ADLIB_INST/GPI[19]INT_NET\, GPI(18) => 
        \Intro_0/MSS_ADLIB_INST/GPI[18]INT_NET\, GPI(17) => 
        \Intro_0/MSS_ADLIB_INST/GPI[17]INT_NET\, GPI(16) => 
        \Intro_0/MSS_ADLIB_INST/GPI[16]INT_NET\, GPI(15) => 
        GLMUXINT_GND, GPI(14) => GLMUXINT_GND, GPI(13) => 
        GLMUXINT_GND, GPI(12) => GLMUXINT_GND, GPI(11) => 
        GLMUXINT_GND, GPI(10) => GLMUXINT_GND, GPI(9) => 
        GLMUXINT_GND, GPI(8) => GLMUXINT_GND, GPI(7) => 
        GLMUXINT_GND, GPI(6) => GLMUXINT_GND, GPI(5) => 
        GLMUXINT_GND, GPI(4) => GLMUXINT_GND, GPI(3) => 
        GLMUXINT_GND, GPI(2) => GLMUXINT_GND, GPI(1) => 
        GLMUXINT_GND, GPI(0) => GLMUXINT_GND, GPO(31) => 
        \Intro_0/MSS_ADLIB_INST/GPO[31]INT_NET\, GPO(30) => 
        \Intro_0/MSS_ADLIB_INST/GPO[30]INT_NET\, GPO(29) => 
        \Intro_0/MSS_ADLIB_INST/GPO[29]INT_NET\, GPO(28) => 
        \Intro_0/MSS_ADLIB_INST/GPO[28]INT_NET\, GPO(27) => 
        \Intro_0/MSS_ADLIB_INST/GPO[27]INT_NET\, GPO(26) => 
        \Intro_0/MSS_ADLIB_INST/GPO[26]INT_NET\, GPO(25) => 
        \Intro_0/MSS_ADLIB_INST/GPO[25]INT_NET\, GPO(24) => 
        \Intro_0/MSS_ADLIB_INST/GPO[24]INT_NET\, GPO(23) => 
        \Intro_0/MSS_ADLIB_INST/GPO[23]INT_NET\, GPO(22) => 
        \Intro_0/MSS_ADLIB_INST/GPO[22]INT_NET\, GPO(21) => 
        \Intro_0/MSS_ADLIB_INST/GPO[21]INT_NET\, GPO(20) => 
        \Intro_0/MSS_ADLIB_INST/GPO[20]INT_NET\, GPO(19) => 
        \Intro_0/MSS_ADLIB_INST/GPO[19]INT_NET\, GPO(18) => 
        \Intro_0/MSS_ADLIB_INST/GPO[18]INT_NET\, GPO(17) => 
        \Intro_0/MSS_ADLIB_INST/GPO[17]INT_NET\, GPO(16) => 
        \Intro_0/MSS_ADLIB_INST/GPO[16]INT_NET\, GPO(15) => nc88, 
        GPO(14) => nc53, GPO(13) => nc39, GPO(12) => nc8, GPO(11)
         => nc82, GPO(10) => nc81, GPO(9) => nc79, GPO(8) => nc43, 
        GPO(7) => nc69, GPO(6) => nc56, GPO(5) => nc20, GPO(4)
         => nc10, GPO(3) => nc57, GPO(2) => nc95, GPO(1) => nc24, 
        GPO(0) => nc14, MACM2FTXD(1) => nc46, MACM2FTXD(0) => 
        nc30, MACF2MRXD(1) => GLMUXINT_GND, MACF2MRXD(0) => 
        GLMUXINT_GND, ACEFLAGS(31) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[31]INT_NET\, 
        ACEFLAGS(30) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[30]INT_NET\, 
        ACEFLAGS(29) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[29]INT_NET\, 
        ACEFLAGS(28) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[28]INT_NET\, 
        ACEFLAGS(27) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[27]INT_NET\, 
        ACEFLAGS(26) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[26]INT_NET\, 
        ACEFLAGS(25) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[25]INT_NET\, 
        ACEFLAGS(24) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[24]INT_NET\, 
        ACEFLAGS(23) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[23]INT_NET\, 
        ACEFLAGS(22) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[22]INT_NET\, 
        ACEFLAGS(21) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[21]INT_NET\, 
        ACEFLAGS(20) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[20]INT_NET\, 
        ACEFLAGS(19) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[19]INT_NET\, 
        ACEFLAGS(18) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[18]INT_NET\, 
        ACEFLAGS(17) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[17]INT_NET\, 
        ACEFLAGS(16) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[16]INT_NET\, 
        ACEFLAGS(15) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[15]INT_NET\, 
        ACEFLAGS(14) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[14]INT_NET\, 
        ACEFLAGS(13) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[13]INT_NET\, 
        ACEFLAGS(12) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[12]INT_NET\, 
        ACEFLAGS(11) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[11]INT_NET\, 
        ACEFLAGS(10) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[10]INT_NET\, ACEFLAGS(9)
         => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[9]INT_NET\, 
        ACEFLAGS(8) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[8]INT_NET\, ACEFLAGS(7)
         => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[7]INT_NET\, 
        ACEFLAGS(6) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[6]INT_NET\, ACEFLAGS(5)
         => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[5]INT_NET\, 
        ACEFLAGS(4) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[4]INT_NET\, ACEFLAGS(3)
         => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[3]INT_NET\, 
        ACEFLAGS(2) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[2]INT_NET\, ACEFLAGS(1)
         => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[1]INT_NET\, 
        ACEFLAGS(0) => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[0]INT_NET\, UART0CTSn
         => \Intro_0/MSS_ADLIB_INST/UART0CTSnINT_NET\, UART0DSRn
         => \Intro_0/MSS_ADLIB_INST/UART0DSRnINT_NET\, UART0RTSn
         => \Intro_0/MSS_ADLIB_INST/UART0RTSnINT_NET\, UART0DTRn
         => \Intro_0/MSS_ADLIB_INST/UART0DTRnINT_NET\, UART0RIn
         => \Intro_0/MSS_ADLIB_INST/UART0RInINT_NET\, UART0DCDn
         => \Intro_0/MSS_ADLIB_INST/UART0DCDnINT_NET\, UART1CTSn
         => \Intro_0/MSS_ADLIB_INST/UART1CTSnINT_NET\, UART1DSRn
         => \Intro_0/MSS_ADLIB_INST/UART1DSRnINT_NET\, UART1RIn
         => \Intro_0/MSS_ADLIB_INST/UART1RInINT_NET\, UART1DCDn
         => \Intro_0/MSS_ADLIB_INST/UART1DCDnINT_NET\, 
        I2C0SMBALERTNO => 
        \Intro_0/MSS_ADLIB_INST/I2C0SMBALERTNOINT_NET\, I2C0BCLK
         => \Intro_0/MSS_ADLIB_INST/I2C0BCLKINT_NET\, 
        I2C0SMBALERTNI => 
        \Intro_0/MSS_ADLIB_INST/I2C0SMBALERTNIINT_NET\, 
        I2C0SMBUSNI => 
        \Intro_0/MSS_ADLIB_INST/I2C0SMBUSNIINT_NET\, 
        I2C1SMBALERTNO => 
        \Intro_0/MSS_ADLIB_INST/I2C1SMBALERTNOINT_NET\, I2C1BCLK
         => \Intro_0/MSS_ADLIB_INST/I2C1BCLKINT_NET\, 
        I2C1SMBALERTNI => 
        \Intro_0/MSS_ADLIB_INST/I2C1SMBALERTNIINT_NET\, 
        I2C1SMBUSNI => 
        \Intro_0/MSS_ADLIB_INST/I2C1SMBUSNIINT_NET\, UART1RTSn
         => \Intro_0/MSS_ADLIB_INST/UART1RTSnINT_NET\, UART1DTRn
         => \Intro_0/MSS_ADLIB_INST/UART1DTRnINT_NET\, TXEV => 
        \Intro_0/MSS_ADLIB_INST/TXEVINT_NET\, RXEV => 
        \Intro_0/MSS_ADLIB_INST/RXEVINT_NET\, VRON => 
        \Intro_0/MSS_ADLIB_INST/VRONINT_NET\, MACM2FTXEN => OPEN, 
        MACF2MCRSDV => GLMUXINT_GND, MACM2FMDEN => OPEN, 
        MACF2MRXER => GLMUXINT_GND, MACM2FMDO => OPEN, MACF2MMDI
         => GLMUXINT_GND, MACM2FMDC => OPEN, I2C0SMBUSNO => 
        \Intro_0/MSS_ADLIB_INST/I2C0SMBUSNOINT_NET\, I2C1SMBUSNO
         => \Intro_0/MSS_ADLIB_INST/I2C1SMBUSNOINT_NET\, CALIBOUT
         => \Intro_0/MSS_ADLIB_INST/CALIBOUTINT_NET\, CALIBIN => 
        \Intro_0/MSS_ADLIB_INST/CALIBININT_NET\, LVTTL0 => 
        \Intro_0/MSS_ADLIB_INST/LVTTL0INT_NET\, LVTTL1 => 
        \Intro_0/MSS_ADLIB_INST/LVTTL1INT_NET\, LVTTL2 => 
        \Intro_0/MSS_ADLIB_INST/LVTTL2INT_NET\, LVTTL0EN => 
        \Intro_0/MSS_ADLIB_INST/LVTTL0ENINT_NET\, LVTTL1EN => 
        \Intro_0/MSS_ADLIB_INST/LVTTL1ENINT_NET\, LVTTL2EN => 
        \Intro_0/MSS_ADLIB_INST/LVTTL2ENINT_NET\, LVTTL3 => 
        \Intro_0/MSS_ADLIB_INST/LVTTL3INT_NET\, LVTTL4 => 
        \Intro_0/MSS_ADLIB_INST/LVTTL4INT_NET\, LVTTL5 => 
        \Intro_0/MSS_ADLIB_INST/LVTTL5INT_NET\, LVTTL3EN => 
        \Intro_0/MSS_ADLIB_INST/LVTTL3ENINT_NET\, LVTTL4EN => 
        \Intro_0/MSS_ADLIB_INST/LVTTL4ENINT_NET\, LVTTL5EN => 
        \Intro_0/MSS_ADLIB_INST/LVTTL5ENINT_NET\, LVTTL6 => 
        \Intro_0/MSS_ADLIB_INST/LVTTL6INT_NET\, LVTTL7 => 
        \Intro_0/MSS_ADLIB_INST/LVTTL7INT_NET\, LVTTL8 => OPEN, 
        LVTTL6EN => \Intro_0/MSS_ADLIB_INST/LVTTL6ENINT_NET\, 
        LVTTL7EN => \Intro_0/MSS_ADLIB_INST/LVTTL7ENINT_NET\, 
        LVTTL8EN => OPEN, LVTTL9 => OPEN, LVTTL10 => OPEN, 
        LVTTL11 => OPEN, LVTTL9EN => OPEN, LVTTL10EN => OPEN, 
        LVTTL11EN => OPEN, CMP0 => 
        \Intro_0/MSS_ADLIB_INST/CMP0INT_NET\, CMP1 => 
        \Intro_0/MSS_ADLIB_INST/CMP1INT_NET\, CMP2 => 
        \Intro_0/MSS_ADLIB_INST/CMP2INT_NET\, CMP3 => 
        \Intro_0/MSS_ADLIB_INST/CMP3INT_NET\, CMP4 => 
        \Intro_0/MSS_ADLIB_INST/CMP4INT_NET\, CMP5 => 
        \Intro_0/MSS_ADLIB_INST/CMP5INT_NET\, FABSDD0D => 
        \Intro_0/MSS_ADLIB_INST/FABSDD0DINT_NET\, FABSDD1D => 
        \Intro_0/MSS_ADLIB_INST/FABSDD1DINT_NET\, FABSDD2D => 
        OPEN, CMP6 => \Intro_0/MSS_ADLIB_INST/CMP6INT_NET\, CMP7
         => \Intro_0/MSS_ADLIB_INST/CMP7INT_NET\, CMP8 => OPEN, 
        FABACETRIG => \Intro_0/MSS_ADLIB_INST/FABACETRIGINT_NET\, 
        CMP9 => OPEN, FABSDD0CLK => 
        \Intro_0/MSS_ADLIB_INST/FABSDD0CLKINT_NET\, FABSDD1CLK
         => \Intro_0/MSS_ADLIB_INST/FABSDD1CLKINT_NET\, 
        FABSDD2CLK => OPEN, VCC15GOOD => 
        \Intro_0/MSS_ADLIB_INST/VCC15GOODINT_NET\, VCC33GOOD => 
        \Intro_0/MSS_ADLIB_INST/VCC33GOODINT_NET\, PUFABn => 
        \Intro_0/MSS_ADLIB_INST/PUFABnINT_NET\, MSSPREADY => 
        \Intro_0/MSS_ADLIB_INST/MSSPREADYINT_NET\, MSSPSLVERR => 
        \Intro_0/MSS_ADLIB_INST/MSSPSLVERRINT_NET\, MSSPSEL => 
        \Intro_0/MSS_ADLIB_INST/MSSPSELINT_NET\, MSSPENABLE => 
        \Intro_0/MSS_ADLIB_INST/MSSPENABLEINT_NET\, MSSPWRITE => 
        \Intro_0/MSS_ADLIB_INST/MSSPWRITEINT_NET\, FABPSEL => 
        \Intro_0/MSS_ADLIB_INST/FABPSELINT_NET\, FABPENABLE => 
        \Intro_0/MSS_ADLIB_INST/FABPENABLEINT_NET\, FABPWRITE => 
        \Intro_0/MSS_ADLIB_INST/FABPWRITEINT_NET\, FABPREADY => 
        \Intro_0/MSS_ADLIB_INST/FABPREADYINT_NET\, FABPSLVERR => 
        \Intro_0/MSS_ADLIB_INST/FABPSLVERRINT_NET\, DEEPSLEEP => 
        \Intro_0/MSS_ADLIB_INST/DEEPSLEEPINT_NET\, SLEEP => 
        \Intro_0/MSS_ADLIB_INST/SLEEPINT_NET\, M2FRESETn => 
        \Intro_0/MSS_ADLIB_INST/M2FRESETnINT_NET\, WDINT => 
        \Intro_0/MSS_ADLIB_INST/WDINTINT_NET\, FABINT => 
        \Intro_0/MSS_ADLIB_INST/FABINTINT_NET\, F2MRESETn => 
        \Intro_0/MSS_ADLIB_INST/F2MRESETnINT_NET\, SYNCCLKFDBK
         => \Intro_0/MSS_ADLIB_INST/SYNCCLKFDBKINT_NET\, CMP10
         => OPEN, CMP11 => OPEN);
    
    \FlashLED_control_wrapper_0/M1/REG_control[4]\ : DLN1
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[4]\, G => 
        \FlashLED_control_wrapper_0/M1/REG_control_0_sqmuxa_net_1\, 
        Q => \FlashLED_control_wrapper_0/M1/REG_control[4]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO_0[13]\ : NOR2B
      port map(A => \CoreTimer_0/DataOut_0_sqmuxa\, B => 
        \CoreTimer_0/Load[13]_net_1\, Y => 
        \CoreTimer_0/Load_m[13]\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_29\ : NOR3C
      port map(A => \CoreAPB3_0.iPSELS_raw_0[1]\, B => 
        \CoreAPB3_0.iPSELS_raw_1[1]\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[29]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[29]\);
    
    \CoreTimer_0/Count[10]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[10]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte_0\, Q => 
        \CoreTimer_0/Count[10]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_55\ : MSS_IF
      port map(PIN4 => \Intro_0_MSS_MASTER_APB_PRDATA[23]\, PIN5
         => \Intro_0_MSS_MASTER_APB_PRDATA[22]\, PIN6 => 
        \Intro_0_MSS_MASTER_APB_PRDATA[24]\, PIN1 => 
        \CoreAPB3_0_APBmslave0_PWDATA[22]\, PIN2 => 
        \CoreAPB3_0_APBmslave0_PWDATA[23]\, PIN3 => 
        \CoreAPB3_0_APBmslave0_PWDATA[24]\, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[23]INT_NET\, PIN5INT
         => \Intro_0/MSS_ADLIB_INST/MSSPRDATA[22]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/MSSPRDATA[24]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[22]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[23]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[24]INT_NET\);
    
    \CoreTimer_0/iPRDATA_RNO_0[20]\ : MX2
      port map(A => \CoreTimer_0/Load[20]_net_1\, B => 
        \CoreTimer_0/Count[20]_net_1\, S => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, Y => 
        \CoreTimer_0/iPRDATA_RNO_0[20]_net_1\);
    
    \CoreTimer_0/Count_RNI29BK1[4]\ : OR2
      port map(A => \CoreTimer_0/Count_c3\, B => 
        \CoreTimer_0/Count[4]_net_1\, Y => \CoreTimer_0/Count_c4\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_13\ : NOR3C
      port map(A => \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, B => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[13]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[13]\);
    
    \CoreTimer_0/iPRDATA_RNO_0[9]\ : NOR2B
      port map(A => \CoreTimer_0/DataOut_0_sqmuxa\, B => 
        \CoreTimer_0/Load[9]_net_1\, Y => \CoreTimer_0/Load_m[9]\);
    
    \FlashLED_control_wrapper_0/M1/REG_load_value[4]\ : DLN1
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[4]\, G => 
        \FlashLED_control_wrapper_0/M1/REG_control_1_sqmuxa_net_1\, 
        Q => 
        \FlashLED_control_wrapper_0/M1/REG_load_value[4]_net_1\);
    
    \CoreTimer_0/Load[31]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[31]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\, Q => 
        \CoreTimer_0/Load[31]_net_1\);
    
    \Intro_0/MSS_SPI_0_SS\ : IOPAD_BI
      port map(D => \Intro_0/SPI0SSO_net_0[0]\, E => 
        \Intro_0/MSS_SPI_0_SS_E\, Y => \Intro_0/MSS_SPI_0_SS_Y\, 
        PAD => SPI_0_SS);
    
    \CoreTimer_0/PreScale_RNIIAR5[8]\ : OR3A
      port map(A => \CoreTimer_0/PreScale[7]_net_1\, B => 
        \CoreTimer_0/N_152\, C => \CoreTimer_0/PreScale_i_0[8]\, 
        Y => \CoreTimer_0/N_441\);
    
    \CoreTimer_0/Count[25]\ : DFN1E1P0
      port map(D => \CoreTimer_0/N_392\, CLK => FAB_CLK, PRE => 
        Intro_0_M2F_RESET_N, E => \CoreTimer_0/Counte_0\, Q => 
        \CoreTimer_0/Count[25]_net_1\);
    
    \FlashLED_control_wrapper_0/M1/RD[4]\ : DLN1
      port map(D => 
        \FlashLED_control_wrapper_0/M1/REG_load_value[4]_net_1\, 
        G => \FlashLED_control_wrapper_0/M1/un2_rwclk\, Q => 
        \RD_c[4]\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_23\ : NOR3C
      port map(A => \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, B => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[23]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[23]\);
    
    \CoreTimer_0/iPRDATA_RNO[9]\ : AO1
      port map(A => \CoreTimer_0/DataOut_1_sqmuxa\, B => 
        \CoreTimer_0/Count[9]_net_1\, C => 
        \CoreTimer_0/Load_m[9]\, Y => \CoreTimer_0/PrdataNext[9]\);
    
    \CoreTimer_0/iPRDATA_RNO[22]\ : NOR3A
      port map(A => \CoreTimer_0/iPRDATA_RNO_0[22]_net_1\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, C => 
        \CoreTimer_0/N_151\, Y => \CoreTimer_0/N_119\);
    
    \CoreTimer_0/Count[2]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[2]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte\, Q => \CoreTimer_0/Count[2]_net_1\);
    
    \CoreTimer_0/Count[28]\ : DFN1E1P0
      port map(D => \CoreTimer_0/N_395\, CLK => FAB_CLK, PRE => 
        Intro_0_M2F_RESET_N, E => \CoreTimer_0/Counte\, Q => 
        \CoreTimer_0/Count[28]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO_0[31]\ : NOR2B
      port map(A => \CoreTimer_0/DataOut_0_sqmuxa\, B => 
        \CoreTimer_0/Load[31]_net_1\, Y => 
        \CoreTimer_0/Load_m[31]\);
    
    \CoreTimer_0/Count_RNO[5]\ : AX1B
      port map(A => \CoreTimer_0/Count_c4\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_184\, Y
         => \CoreTimer_0/Count_RNO[5]_net_1\);
    
    \RD_pad[7]/U0/U1\ : IOTRI_OB_EB
      port map(D => \RD_c[7]\, E => PLLEN_VCC, DOUT => 
        \RD_pad[7]/U0/NET1\, EOUT => \RD_pad[7]/U0/NET2\);
    
    \CoreTimer_0/Load[0]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[0]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0\, Q => 
        \CoreTimer_0/Load[0]_net_1\);
    
    \RD_pad[4]/U0/U0\ : IOPAD_TRI
      port map(D => \RD_pad[4]/U0/NET1\, E => \RD_pad[4]/U0/NET2\, 
        PAD => RD(4));
    
    \CoreTimer_0/Count_RNO[31]\ : AX1B
      port map(A => \CoreTimer_0/Count_c29\, B => 
        \CoreTimer_0/Count_66_0\, C => \CoreTimer_0/N_236\, Y => 
        \CoreTimer_0/Count_RNO[31]_net_1\);
    
    \CoreTimer_0/TimerPre[2]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[2]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_prescaleen_0_a2_1_a3_net_1\, Q => 
        \CoreTimer_0/TimerPre[2]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO_1[2]\ : NOR3B
      port map(A => \CoreAPB3_0_APBmslave0_PADDR_0[3]\, B => 
        \CoreAPB3_0_APBmslave0_PADDR_0[2]\, C => 
        \CoreTimer_0/TimerPre[2]_net_1\, Y => \CoreTimer_0/N_239\);
    
    \CoreTimer_0/Count_RNIB2DV[2]\ : OR2
      port map(A => \CoreTimer_0/N_153\, B => 
        \CoreTimer_0/Count[2]_net_1\, Y => \CoreTimer_0/N_154\);
    
    \CoreTimer_0/Load[15]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[15]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0\, Q => 
        \CoreTimer_0/Load[15]_net_1\);
    
    \CoreTimer_0/Load[2]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[2]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0\, Q => 
        \CoreTimer_0/Load[2]_net_1\);
    
    \CoreTimer_0/Load[20]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[20]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\, Q => 
        \CoreTimer_0/Load[20]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO[6]\ : AO1
      port map(A => \CoreTimer_0/DataOut_1_sqmuxa\, B => 
        \CoreTimer_0/Count[6]_net_1\, C => 
        \CoreTimer_0/Load_m[6]\, Y => \CoreTimer_0/PrdataNext[6]\);
    
    \Intro_0/MSS_ADLIB_INST/U_90\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[29]INT_NET\, PIN5INT
         => \Intro_0/MSS_ADLIB_INST/FABPWDATA[28]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/FABPWDATA[30]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[28]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[29]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[30]INT_NET\);
    
    \CoreTimer_0/iPRDATA_RNO[25]\ : AO1
      port map(A => \CoreTimer_0/DataOut_1_sqmuxa\, B => 
        \CoreTimer_0/Count[25]_net_1\, C => 
        \CoreTimer_0/Load_m[25]\, Y => 
        \CoreTimer_0/PrdataNext[25]\);
    
    \CoreTimer_0/iPRDATA[5]\ : DFN1C0
      port map(D => \CoreTimer_0/PrdataNext[5]\, CLK => FAB_CLK, 
        CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[5]\);
    
    \CoreTimer_0/Count_RNIRKU51[28]\ : OR3
      port map(A => \CoreTimer_0/Count[28]_net_1\, B => 
        \CoreTimer_0/Count[29]_net_1\, C => 
        \CoreTimer_0/N_58_i_0_o2_12\, Y => 
        \CoreTimer_0/N_58_i_0_o2_20\);
    
    \CoreTimer_0/Count[0]\ : DFN1P0
      port map(D => \CoreTimer_0/N_507_mux\, CLK => FAB_CLK, PRE
         => Intro_0_M2F_RESET_N, Q => 
        \CoreTimer_0/Count[0]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_88\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[23]INT_NET\, PIN5INT
         => \Intro_0/MSS_ADLIB_INST/FABPWDATA[22]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/FABPWDATA[24]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[22]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[23]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[24]INT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_48\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[2]INT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[1]INT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[3]INT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[1]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[2]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[3]INT_NET\);
    
    \CoreTimer_0/Count_RNIKTVN4[14]\ : OR2
      port map(A => \CoreTimer_0/Count_c13\, B => 
        \CoreTimer_0/Count[14]_net_1\, Y => 
        \CoreTimer_0/Count_c14\);
    
    \CoreAPB3_0/iPSELS_raw_0[1]\ : NOR3A
      port map(A => Intro_0_MSS_MASTER_APB_PSELx, B => 
        \Intro_0_MSS_MASTER_APB_PADDR[11]\, C => 
        \Intro_0_MSS_MASTER_APB_PADDR[10]\, Y => 
        \CoreAPB3_0.iPSELS_raw_0[1]\);
    
    \Intro_0/MSS_ADLIB_INST/U_62\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => \Intro_0/MSS_ADLIB_INST/LVTTL1ENINT_NET\, 
        PIN5INT => \Intro_0/MSS_ADLIB_INST/LVTTL0ENINT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/LVTTL2ENINT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/LVTTL0INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/LVTTL1INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/LVTTL2INT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_6\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => \Intro_0/MSS_ADLIB_INST/GPI[29]INT_NET\, 
        PIN5INT => \Intro_0/MSS_ADLIB_INST/GPI[28]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/GPI[30]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/GPO[28]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/GPO[29]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/GPO[30]INT_NET\);
    
    \CoreTimer_0/iPRDATA_RNO_0[18]\ : MX2
      port map(A => \CoreTimer_0/Load[18]_net_1\, B => 
        \CoreTimer_0/Count[18]_net_1\, S => 
        \CoreAPB3_0_APBmslave0_PADDR_0[2]\, Y => 
        \CoreTimer_0/N_455\);
    
    \FlashLED_control_wrapper_0/M1/RD[7]\ : DLN1
      port map(D => 
        \FlashLED_control_wrapper_0/M1/REG_load_value[7]_net_1\, 
        G => \FlashLED_control_wrapper_0/M1/un2_rwclk\, Q => 
        \RD_c[7]\);
    
    \FlashLED_control_wrapper_0/M1/RD[6]\ : DLN1
      port map(D => 
        \FlashLED_control_wrapper_0/M1/REG_load_value[6]_net_1\, 
        G => \FlashLED_control_wrapper_0/M1/un2_rwclk\, Q => 
        \RD_c[6]\);
    
    \CoreTimer_0/Count[14]\ : DFN1E1P0
      port map(D => \CoreTimer_0/N_381\, CLK => FAB_CLK, PRE => 
        Intro_0_M2F_RESET_N, E => \CoreTimer_0/Counte_0\, Q => 
        \CoreTimer_0/Count[14]_net_1\);
    
    \CoreTimer_0/Count[4]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[4]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte\, Q => \CoreTimer_0/Count[4]_net_1\);
    
    \CoreTimer_0/Count_RNO[1]\ : MX2A
      port map(A => \CoreTimer_0/N_190_i\, B => 
        \CoreTimer_0/Load[1]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => 
        \CoreTimer_0/Count_RNO[1]_net_1\);
    
    \CoreTimer_0/CountPulse_RNO_3\ : NOR2
      port map(A => \CoreTimer_0/TimerPre[1]_net_1\, B => 
        \CoreTimer_0/TimerPre[2]_net_1\, Y => 
        \CoreTimer_0/NextCountPulse_0_0_a3_4_0\);
    
    \Intro_0/MSS_SPI_0_DI\ : IOPAD_IN
      port map(PAD => SPI_0_DI, Y => \Intro_0/MSS_SPI_0_DI_Y\);
    
    \CoreTimer_0/iPRDATA[2]\ : DFN1C0
      port map(D => \CoreTimer_0/iPRDATA_RNO[2]_net_1\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[2]\);
    
    \CoreTimer_0/Count_RNINMS91[4]\ : OR3
      port map(A => \CoreTimer_0/Count[4]_net_1\, B => 
        \CoreTimer_0/Count[8]_net_1\, C => 
        \CoreTimer_0/N_58_i_0_o2_4\, Y => 
        \CoreTimer_0/N_58_i_0_o2_16\);
    
    \CoreTimer_0/Count_RNIG9KR3[11]\ : OR2
      port map(A => \CoreTimer_0/Count_c10\, B => 
        \CoreTimer_0/Count[11]_net_1\, Y => 
        \CoreTimer_0/Count_c11\);
    
    \Intro_0/MSS_ADLIB_INST/U_2\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => \Intro_0/MSS_ADLIB_INST/GPI[17]INT_NET\, 
        PIN5INT => \Intro_0/MSS_ADLIB_INST/GPI[16]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/GPI[18]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/GPO[16]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/GPO[17]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/GPO[18]INT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_85\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[29]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[30]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[31]INT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_59\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => GLMUXINT_GND, PIN2INT => GLMUXINT_GND, PIN3INT
         => GLMUXINT_GND);
    
    \Intro_0/MSS_ADLIB_INST/U_45\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[25]INT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[24]INT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[26]INT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/MSSINT[2]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/MSSINT[3]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/MSSINT[4]INT_NET\);
    
    \CoreTimer_0/PrdataNext_0_iv_0_i_a2[3]\ : NOR2A
      port map(A => \CoreAPB3_0_APBmslave0_PADDR[3]\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, Y => 
        \CoreTimer_0/N_257\);
    
    \CoreTimer_0/iPRDATA_RNO_7[0]\ : NOR3A
      port map(A => \CoreTimer_0/N_257\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, C => 
        \CoreTimer_0/CtrlReg[0]_net_1\, Y => \CoreTimer_0/N_492\);
    
    \CoreTimer_0/iPRDATA_RNO_0[4]\ : NOR2B
      port map(A => \CoreTimer_0/DataOut_0_sqmuxa\, B => 
        \CoreTimer_0/Load[4]_net_1\, Y => \CoreTimer_0/Load_m[4]\);
    
    \Intro_0/MSS_ADLIB_INST/U_67\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => GLMUXINT_GND, PIN2INT => GLMUXINT_GND, PIN3INT
         => GLMUXINT_GND);
    
    \CoreTimer_0/PreScale[3]\ : DFN1C0
      port map(D => \CoreTimer_0/N_26\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => \CoreTimer_0/PreScale[3]_net_1\);
    
    \CoreTimer_0/Load[4]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[4]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0\, Q => 
        \CoreTimer_0/Load[4]_net_1\);
    
    \CoreTimer_0/Count_RNO[29]\ : AX1B
      port map(A => \CoreTimer_0/un1_loadenreg\, B => 
        \CoreTimer_0/Count_c28\, C => \CoreTimer_0/N_232\, Y => 
        \CoreTimer_0/N_396\);
    
    \CoreTimer_0/Count_RNIRP254[12]\ : OR2
      port map(A => \CoreTimer_0/Count_c11\, B => 
        \CoreTimer_0/Count[12]_net_1\, Y => 
        \CoreTimer_0/Count_c12\);
    
    \CoreTimer_0/iPRDATA_RNO[17]\ : AO1
      port map(A => \CoreTimer_0/DataOut_1_sqmuxa\, B => 
        \CoreTimer_0/Count[17]_net_1\, C => 
        \CoreTimer_0/Load_m[17]\, Y => 
        \CoreTimer_0/PrdataNext[17]\);
    
    \CoreTimer_0/CtrlReg[1]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[1]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un6_ctrlen_0_a2_0_a2_net_1\, Q => 
        \CoreTimer_0/CtrlReg[1]_net_1\);
    
    \CoreTimer_0/PreScale[2]\ : DFN1P0
      port map(D => \CoreTimer_0/N_28\, CLK => FAB_CLK, PRE => 
        Intro_0_M2F_RESET_N, Q => \CoreTimer_0/PreScale_i_0[2]\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_18\ : NOR3C
      port map(A => \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, B => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[18]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[18]\);
    
    \CoreTimer_0/Count_RNIIHQT5[18]\ : OR2
      port map(A => \CoreTimer_0/Count_c17\, B => 
        \CoreTimer_0/Count[18]_net_1\, Y => 
        \CoreTimer_0/Count_c18\);
    
    \CoreTimer_0/Count_RNI65S91[3]\ : OR2
      port map(A => \CoreTimer_0/N_154\, B => 
        \CoreTimer_0/Count[3]_net_1\, Y => \CoreTimer_0/Count_c3\);
    
    \CoreTimer_0/PreScale_RNI0O73[4]\ : OR2
      port map(A => \CoreTimer_0/PreScale_i_0[4]\, B => 
        \CoreTimer_0/N_146\, Y => \CoreTimer_0/N_148\);
    
    \CoreTimer_0/CountPulse_RNO_9\ : OR2A
      port map(A => \CoreTimer_0/TimerPre[0]_net_1\, B => 
        \CoreTimer_0/PreScale[1]_net_1\, Y => \CoreTimer_0/N_440\);
    
    \CoreTimer_0/LoadEnReg_RNIF830L\ : OR3
      port map(A => \CoreTimer_0/N_248\, B => 
        \CoreTimer_0/LoadEnReg_net_1\, C => 
        \CoreTimer_0/CtrlReg_RNIC1I6A[2]_net_1\, Y => 
        \CoreTimer_0/Counte_0\);
    
    \Intro_0/MSS_ADLIB_INST/U_54\ : MSS_IF
      port map(PIN4 => \Intro_0_MSS_MASTER_APB_PRDATA[20]\, PIN5
         => \Intro_0_MSS_MASTER_APB_PRDATA[19]\, PIN6 => 
        \Intro_0_MSS_MASTER_APB_PRDATA[21]\, PIN1 => 
        \CoreAPB3_0_APBmslave0_PWDATA[19]\, PIN2 => 
        \CoreAPB3_0_APBmslave0_PWDATA[20]\, PIN3 => 
        \CoreAPB3_0_APBmslave0_PWDATA[21]\, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[20]INT_NET\, PIN5INT
         => \Intro_0/MSS_ADLIB_INST/MSSPRDATA[19]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/MSSPRDATA[21]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[19]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[20]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[21]INT_NET\);
    
    \CoreTimer_0/PreScale_RNO[7]\ : XA1C
      port map(A => \CoreTimer_0/N_152\, B => 
        \CoreTimer_0/PreScale[7]_net_1\, C => 
        \CoreTimer_0/N_16_2\, Y => \CoreTimer_0/N_18\);
    
    \CoreTimer_0/iPRDATA_RNO[2]\ : NOR3
      port map(A => \CoreTimer_0/PrdataNext_0_iv_0_i_0[2]\, B => 
        \CoreTimer_0/N_239\, C => 
        \CoreTimer_0/PrdataNext_0_iv_0_i_1[2]\, Y => 
        \CoreTimer_0/iPRDATA_RNO[2]_net_1\);
    
    \CoreTimer_0/Count_RNO_0[5]\ : MX2
      port map(A => \CoreTimer_0/Count[5]_net_1\, B => 
        \CoreTimer_0/Load[5]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_184\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_28\ : NOR3C
      port map(A => \CoreAPB3_0.iPSELS_raw_0[1]\, B => 
        \CoreAPB3_0.iPSELS_raw_1[1]\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[28]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[28]\);
    
    \CoreAPB3_0/iPSELS_raw_1[1]\ : NOR2A
      port map(A => \Intro_0_MSS_MASTER_APB_PADDR[8]\, B => 
        \Intro_0_MSS_MASTER_APB_PADDR[9]\, Y => 
        \CoreAPB3_0.iPSELS_raw_1[1]\);
    
    \CoreTimer_0/Count_RNO_0[17]\ : MX2
      port map(A => \CoreTimer_0/Count[17]_net_1\, B => 
        \CoreTimer_0/Load[17]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_208\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_11\ : NOR3C
      port map(A => \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, B => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[11]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[11]\);
    
    \CoreTimer_0/PreScale_RNO[4]\ : OR3A
      port map(A => \CoreTimer_0/N_148\, B => 
        \CoreTimer_0/PreScale_n4_i_0_0\, C => 
        \CoreTimer_0/CtrlReg_RNIC1I6A[2]_net_1\, Y => 
        \CoreTimer_0/N_24\);
    
    \CoreTimer_0/CtrlReg_RNI9LMM[1]\ : NOR2B
      port map(A => \CoreTimer_0/CtrlReg[1]_net_1\, B => 
        \CoreTimer_0/RawTimInt_net_1\, Y => \CoreTimer_0.N_10\);
    
    \CoreAPB3_0/iPSELS_raw_0_0[1]\ : NOR3A
      port map(A => Intro_0_MSS_MASTER_APB_PSELx, B => 
        \Intro_0_MSS_MASTER_APB_PADDR[11]\, C => 
        \Intro_0_MSS_MASTER_APB_PADDR[10]\, Y => 
        \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO_0[29]\ : MX2
      port map(A => \CoreTimer_0/Load[29]_net_1\, B => 
        \CoreTimer_0/Count[29]_net_1\, S => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, Y => 
        \CoreTimer_0/N_461\);
    
    \CoreTimer_0/Count[23]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[23]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte_0\, Q => 
        \CoreTimer_0/Count[23]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_76\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[2]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[3]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[4]INT_NET\);
    
    \CoreTimer_0/Count[29]\ : DFN1E1P0
      port map(D => \CoreTimer_0/N_396\, CLK => FAB_CLK, PRE => 
        Intro_0_M2F_RESET_N, E => \CoreTimer_0/Counte\, Q => 
        \CoreTimer_0/Count[29]_net_1\);
    
    \CoreTimer_0/Count_RNIEPOG6[20]\ : OR2
      port map(A => \CoreTimer_0/Count_c19\, B => 
        \CoreTimer_0/Count[20]_net_1\, Y => 
        \CoreTimer_0/Count_c20\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_21\ : NOR3C
      port map(A => \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, B => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[21]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[21]\);
    
    \Intro_0/MSS_RESET_0_MSS_RESET_N\ : IOPAD_IN
      port map(PAD => MSS_RESET_N, Y => 
        \Intro_0/MSS_RESET_0_MSS_RESET_N_Y\);
    
    \CoreTimer_0/TimerPre[3]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[3]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_prescaleen_0_a2_1_a3_net_1\, Q => 
        \CoreTimer_0/TimerPre[3]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_60\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => \CoreTimer_0.N_10\, 
        PIN6 => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3
         => OPEN, PIN4INT => OPEN, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/FABINTINT_NET\, PIN6INT => OPEN, 
        PIN1INT => GLMUXINT_GND, PIN2INT => GLMUXINT_GND, PIN3INT
         => GLMUXINT_GND);
    
    \CoreTimer_0/iPRDATA_RNO_0[17]\ : NOR2B
      port map(A => \CoreTimer_0/DataOut_0_sqmuxa\, B => 
        \CoreTimer_0/Load[17]_net_1\, Y => 
        \CoreTimer_0/Load_m[17]\);
    
    \Intro_0/MSS_SPI_0_CLK\ : IOPAD_BI
      port map(D => \Intro_0/MSS_SPI_0_CLK_D\, E => 
        \Intro_0/MSS_SPI_0_SS_E\, Y => \Intro_0/MSS_SPI_0_CLK_Y\, 
        PAD => SPI_0_CLK);
    
    \CoreTimer_0/iPRDATA_RNO[19]\ : NOR3A
      port map(A => \CoreTimer_0/iPRDATA_RNO_0[19]_net_1\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, C => 
        \CoreTimer_0/N_151\, Y => \CoreTimer_0/N_113\);
    
    \CoreTimer_0/Count_RNI1EVI[26]\ : OR2
      port map(A => \CoreTimer_0/Count[26]_net_1\, B => 
        \CoreTimer_0/Count[27]_net_1\, Y => 
        \CoreTimer_0/N_58_i_0_o2_1\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_10\ : NOR3C
      port map(A => \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, B => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[10]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[10]\);
    
    \CoreTimer_0/iPRDATA[27]\ : DFN1C0
      port map(D => \CoreTimer_0/PrdataNext[27]\, CLK => FAB_CLK, 
        CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[27]\);
    
    \CoreTimer_0/Count[6]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[6]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte\, Q => \CoreTimer_0/Count[6]_net_1\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_6\ : NOR3C
      port map(A => \CoreAPB3_0.iPSELS_raw_0[1]\, B => 
        \CoreAPB3_0.iPSELS_raw_1[1]\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[6]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[6]\);
    
    \Intro_0/MSS_ADLIB_INST/U_53\ : MSS_IF
      port map(PIN4 => \Intro_0_MSS_MASTER_APB_PRDATA[17]\, PIN5
         => \Intro_0_MSS_MASTER_APB_PRDATA[16]\, PIN6 => 
        \Intro_0_MSS_MASTER_APB_PRDATA[18]\, PIN1 => 
        \CoreAPB3_0_APBmslave0_PWDATA[16]\, PIN2 => 
        \CoreAPB3_0_APBmslave0_PWDATA[17]\, PIN3 => 
        \CoreAPB3_0_APBmslave0_PWDATA[18]\, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[17]INT_NET\, PIN5INT
         => \Intro_0/MSS_ADLIB_INST/MSSPRDATA[16]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/MSSPRDATA[18]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[16]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[17]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[18]INT_NET\);
    
    \FlashLED_control_wrapper_0/M1/REG_control_RNIH4US[6]\ : NOR2
      port map(A => 
        \FlashLED_control_wrapper_0/M1/REG_control[6]_net_1\, B
         => \FlashLED_control_wrapper_0/M1/REG_control[7]_net_1\, 
        Y => \FlashLED_control_wrapper_0/M1/un2_rwclk_3\);
    
    \CoreTimer_0/PreScale[9]\ : DFN1C0
      port map(D => \CoreTimer_0/N_136\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => \CoreTimer_0/PreScale[9]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO[28]\ : NOR3A
      port map(A => \CoreTimer_0/N_460\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, C => 
        \CoreTimer_0/N_151\, Y => \CoreTimer_0/N_121\);
    
    \Intro_0/MSS_ADLIB_INST/U_95\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/I2C1SMBALERTNIINT_NET\, PIN5INT
         => \Intro_0/MSS_ADLIB_INST/I2C1BCLKINT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/I2C1SMBUSNIINT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/SPI1SSO[6]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/SPI1SSO[7]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/I2C1SMBALERTNOINT_NET\);
    
    \CoreTimer_0/Count_RNI49976[19]\ : OR2
      port map(A => \CoreTimer_0/Count_c18\, B => 
        \CoreTimer_0/Count[19]_net_1\, Y => 
        \CoreTimer_0/Count_c19\);
    
    \CoreTimer_0/un5_loaden_0_a2_2_a3_0\ : NOR2B
      port map(A => \CoreTimer_0/N_261\, B => \CoreTimer_0.N_258\, 
        Y => \CoreTimer_0/un5_loaden_0\);
    
    \CoreTimer_0/iPRDATA_RNO_0[6]\ : NOR2B
      port map(A => \CoreTimer_0/DataOut_0_sqmuxa\, B => 
        \CoreTimer_0/Load[6]_net_1\, Y => \CoreTimer_0/Load_m[6]\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_20\ : NOR3C
      port map(A => \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, B => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[20]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[20]\);
    
    \CoreTimer_0/Load[19]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[19]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\, Q => 
        \CoreTimer_0/Load[19]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO[20]\ : NOR3A
      port map(A => \CoreTimer_0/iPRDATA_RNO_0[20]_net_1\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, C => 
        \CoreTimer_0/N_151\, Y => \CoreTimer_0/N_115\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_8\ : NOR3C
      port map(A => \CoreAPB3_0.iPSELS_raw_0[1]\, B => 
        \CoreAPB3_0.iPSELS_raw_1[1]\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[8]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[8]\);
    
    \Intro_0/MSS_ADLIB_INST/U_51\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[11]INT_NET\, PIN5INT
         => \Intro_0/MSS_ADLIB_INST/FABPWDATA[10]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/FABPWDATA[12]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[10]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[11]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[12]INT_NET\);
    
    \FlashLED_control_wrapper_0/M1/REG_control_RNIEKRP1[0]\ : 
        NOR3B
      port map(A => 
        \FlashLED_control_wrapper_0/M1/REG_control[0]_net_1\, B
         => \FlashLED_control_wrapper_0/M1/un2_rwclk_1\, C => 
        \FlashLED_control_wrapper_0/M1/REG_control[1]_net_1\, Y
         => \FlashLED_control_wrapper_0/M1/un2_rwclk_4\);
    
    \CoreTimer_0/Count[12]\ : DFN1E1P0
      port map(D => \CoreTimer_0/N_379\, CLK => FAB_CLK, PRE => 
        Intro_0_M2F_RESET_N, E => \CoreTimer_0/Counte_0\, Q => 
        \CoreTimer_0/Count[12]_net_1\);
    
    \CoreTimer_0/Count_RNI7TPE2[10]\ : OR3
      port map(A => \CoreTimer_0/N_58_i_0_o2_14\, B => 
        \CoreTimer_0/N_58_i_0_o2_13\, C => \CoreTimer_0/N_154\, Y
         => \CoreTimer_0/N_58_i_0_o2_25\);
    
    \Intro_0/MSS_ADLIB_INST/U_89\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[26]INT_NET\, PIN5INT
         => \Intro_0/MSS_ADLIB_INST/FABPWDATA[25]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/FABPWDATA[27]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[25]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[26]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[27]INT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_49\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[5]INT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[4]INT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[6]INT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[4]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[5]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[6]INT_NET\);
    
    \CoreTimer_0/iPRDATA_RNO_0[24]\ : NOR2B
      port map(A => \CoreTimer_0/DataOut_1_sqmuxa\, B => 
        \CoreTimer_0/Count[24]_net_1\, Y => 
        \CoreTimer_0/Count_m[24]\);
    
    \CoreTimer_0/Count[27]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[27]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte\, Q => \CoreTimer_0/Count[27]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO[8]\ : NOR3A
      port map(A => \CoreTimer_0/iPRDATA_RNO_0[8]_net_1\, B => 
        \CoreAPB3_0_APBmslave0_PADDR_0[3]\, C => 
        \CoreTimer_0/N_151\, Y => \CoreTimer_0/N_37\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_15\ : NOR3C
      port map(A => \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, B => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[15]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[15]\);
    
    \CoreTimer_0/Load[27]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[27]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\, Q => 
        \CoreTimer_0/Load[27]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO_8[0]\ : NOR3B
      port map(A => \CoreAPB3_0_APBmslave0_PADDR[4]\, B => 
        \CoreTimer_0/N_448\, C => 
        \CoreAPB3_0_APBmslave0_PADDR_0[2]\, Y => 
        \CoreTimer_0/N_485\);
    
    \CoreTimer_0/iPRDATA[9]\ : DFN1C0
      port map(D => \CoreTimer_0/PrdataNext[9]\, CLK => FAB_CLK, 
        CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[9]\);
    
    \CoreTimer_0/Count_RNIVGM98[26]\ : OR2
      port map(A => \CoreTimer_0/Count_c25\, B => 
        \CoreTimer_0/Count[26]_net_1\, Y => 
        \CoreTimer_0/Count_c26\);
    
    \FlashLED_control_wrapper_0/M1/REG_load_value[0]\ : DLN1
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[0]\, G => 
        \FlashLED_control_wrapper_0/M1/REG_control_1_sqmuxa_net_1\, 
        Q => 
        \FlashLED_control_wrapper_0/M1/REG_load_value[0]_net_1\);
    
    \Intro_0/MSS_UART_0_TXD\ : IOPAD_TRI
      port map(D => \Intro_0/MSS_UART_0_TXD_D\, E => PLLEN_VCC, 
        PAD => UART_0_TXD);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_25\ : NOR3C
      port map(A => \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, B => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[25]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[25]\);
    
    \CoreTimer_0/iPRDATA_RNO_3[3]\ : NOR2
      port map(A => \CoreAPB3_0_APBmslave0_PADDR[2]\, B => 
        \CoreTimer_0/Load[3]_net_1\, Y => \CoreTimer_0/N_244\);
    
    \Intro_0/MSS_ADLIB_INST/U_84\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[26]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[27]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[28]INT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_44\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[22]INT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[21]INT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[23]INT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/SLEEPINT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/MSSINT[0]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/MSSINT[1]INT_NET\);
    
    \CoreTimer_0/Count_RNO_0[10]\ : MX2
      port map(A => \CoreTimer_0/Count[10]_net_1\, B => 
        \CoreTimer_0/Load[10]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_194\);
    
    \CoreTimer_0/Count[3]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[3]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte\, Q => \CoreTimer_0/Count[3]_net_1\);
    
    \CoreTimer_0/Count_RNIN3VI[13]\ : OR2
      port map(A => \CoreTimer_0/Count[30]_net_1\, B => 
        \CoreTimer_0/Count[13]_net_1\, Y => 
        \CoreTimer_0/N_58_i_0_o2_6\);
    
    \CoreTimer_0/Count_RNO[21]\ : AX1B
      port map(A => \CoreTimer_0/Count_c20\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_216\, Y
         => \CoreTimer_0/Count_RNO[21]_net_1\);
    
    \CoreTimer_0/iPRDATA[1]\ : DFN1C0
      port map(D => \CoreTimer_0/N_29\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[1]\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_4\ : NOR3C
      port map(A => \CoreAPB3_0.iPSELS_raw_0[1]\, B => 
        \CoreAPB3_0.iPSELS_raw_1[1]\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[4]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[4]\);
    
    \FlashLED_control_wrapper_0/M1/Write_REGs.un2_wen_1\ : NOR2B
      port map(A => Intro_0_MSS_MASTER_APB_PSELx, B => 
        CoreAPB3_0_APBmslave0_PWRITE, Y => 
        \FlashLED_control_wrapper_0/M1/un2_wen_1\);
    
    \CoreTimer_0/PreScale_RNO[5]\ : NOR3A
      port map(A => \CoreTimer_0/N_150\, B => 
        \CoreTimer_0/PreScale_n5_i_0_0\, C => 
        \CoreTimer_0/CtrlReg_RNIC1I6A[2]_net_1\, Y => 
        \CoreTimer_0/N_22\);
    
    \CoreTimer_0/Count[26]\ : DFN1E1P0
      port map(D => \CoreTimer_0/N_393\, CLK => FAB_CLK, PRE => 
        Intro_0_M2F_RESET_N, E => \CoreTimer_0/Counte_0\, Q => 
        \CoreTimer_0/Count[26]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO_1[0]\ : AO1A
      port map(A => \CoreTimer_0/Count[0]_net_1\, B => 
        \CoreTimer_0/PrdataNext_iv_0_i_a3_3_0[0]\, C => 
        \CoreTimer_0/PrdataNext_iv_0_i_1[0]\, Y => 
        \CoreTimer_0/PrdataNext_iv_0_i_3[0]\);
    
    \FlashLED_control_wrapper_0/M1/REG_control_RNIU4SP1[4]\ : 
        NOR3A
      port map(A => \FlashLED_control_wrapper_0/M1/un2_rwclk_3\, 
        B => \FlashLED_control_wrapper_0/M1/REG_control[5]_net_1\, 
        C => \FlashLED_control_wrapper_0/M1/REG_control[4]_net_1\, 
        Y => \FlashLED_control_wrapper_0/M1/un2_rwclk_5\);
    
    \CoreTimer_0/Count_RNI6Q5I3[10]\ : OR2
      port map(A => \CoreTimer_0/Count_c9\, B => 
        \CoreTimer_0/Count[10]_net_1\, Y => 
        \CoreTimer_0/Count_c10\);
    
    \Intro_0/MSS_ADLIB_INST/U_36\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => PLLEN_VCC, PIN6 => 
        \Intro_0_MSS_MASTER_APB_PRDATA[0]\, PIN1 => OPEN, PIN2
         => OPEN, PIN3 => \CoreAPB3_0_APBmslave0_PWDATA[0]\, 
        PIN4INT => \Intro_0/MSS_ADLIB_INST/MSSPSLVERRINT_NET\, 
        PIN5INT => \Intro_0/MSS_ADLIB_INST/MSSPREADYINT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/MSSPRDATA[0]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/MSSPADDR[18]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/MSSPADDR[19]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[0]INT_NET\);
    
    \CoreTimer_0/IntClr_RNO\ : OR3C
      port map(A => CoreAPB3_0_APBmslave0_PWRITE, B => 
        \CoreTimer_0/N_102\, C => 
        \CoreTimer_0/un5_intclren_0_a3_0_a3_1\, Y => 
        \CoreTimer_0/IntClr_RNO_net_1\);
    
    \CoreTimer_0/Count_RNO_0[2]\ : MX2
      port map(A => \CoreTimer_0/Count[2]_net_1\, B => 
        \CoreTimer_0/Load[2]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_178\);
    
    \CoreTimer_0/Count_RNO[7]\ : AX1B
      port map(A => \CoreTimer_0/Count_c6\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_188\, Y
         => \CoreTimer_0/Count_RNO[7]_net_1\);
    
    \CoreTimer_0/Count_RNO_0[7]\ : MX2
      port map(A => \CoreTimer_0/Count[7]_net_1\, B => 
        \CoreTimer_0/Load[7]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_188\);
    
    \CoreTimer_0/Count_RNO[27]\ : AX1B
      port map(A => \CoreTimer_0/Count_c26\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_228\, Y
         => \CoreTimer_0/Count_RNO[27]_net_1\);
    
    \CoreTimer_0/Count_RNO[26]\ : AX1B
      port map(A => \CoreTimer_0/un1_loadenreg\, B => 
        \CoreTimer_0/Count_c25\, C => \CoreTimer_0/N_226\, Y => 
        \CoreTimer_0/N_393\);
    
    \CoreTimer_0/PreScale[6]\ : DFN1P0
      port map(D => \CoreTimer_0/N_20\, CLK => FAB_CLK, PRE => 
        Intro_0_M2F_RESET_N, Q => \CoreTimer_0/PreScale_i_0[6]\);
    
    \CoreTimer_0/Count_RNO_0[6]\ : MX2
      port map(A => \CoreTimer_0/Count[6]_net_1\, B => 
        \CoreTimer_0/Load[6]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_186\);
    
    \CoreTimer_0/Count[30]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[30]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte\, Q => \CoreTimer_0/Count[30]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_65\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/PUFABnINT_NET\, 
        PIN2INT => GLMUXINT_GND, PIN3INT => GLMUXINT_GND);
    
    \CoreTimer_0/Load[23]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[23]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\, Q => 
        \CoreTimer_0/Load[23]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_83\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[23]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[24]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[25]INT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_43\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[19]INT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[18]INT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[20]INT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/FABPREADYINT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/FABPSLVERRINT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/DEEPSLEEPINT_NET\);
    
    \CoreTimer_0/iPRDATA_RNO_9[0]\ : NOR2A
      port map(A => \CoreTimer_0.N_258\, B => 
        \CoreTimer_0/Load[0]_net_1\, Y => \CoreTimer_0/N_489\);
    
    \CoreTimer_0/Count_RNO_0[13]\ : MX2
      port map(A => \CoreTimer_0/Count[13]_net_1\, B => 
        \CoreTimer_0/Load[13]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_200\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_14\ : NOR3C
      port map(A => \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, B => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[14]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[14]\);
    
    \CoreTimer_0/iPRDATA_RNO_0[8]\ : MX2
      port map(A => \CoreTimer_0/Load[8]_net_1\, B => 
        \CoreTimer_0/Count[8]_net_1\, S => 
        \CoreAPB3_0_APBmslave0_PADDR_0[2]\, Y => 
        \CoreTimer_0/iPRDATA_RNO_0[8]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO_0[2]\ : AO1A
      port map(A => \CoreTimer_0/CtrlReg[2]_net_1\, B => 
        \CoreTimer_0/N_257\, C => \CoreTimer_0/N_151\, Y => 
        \CoreTimer_0/PrdataNext_0_iv_0_i_0[2]\);
    
    \FlashLED_control_wrapper_0/M1/Write_REGs.un2_wen_3\ : NOR3B
      port map(A => \FlashLED_control_wrapper_0/M1/un2_wen_0\, B
         => \FlashLED_control_wrapper_0/M1/un2_wen_1\, C => 
        \Intro_0_MSS_MASTER_APB_PADDR[9]\, Y => 
        \FlashLED_control_wrapper_0/M1/un2_wen_3\);
    
    \CoreTimer_0/DataOut_1_sqmuxa_0_a2_1_a3\ : NOR3A
      port map(A => \CoreAPB3_0_APBmslave0_PADDR[2]\, B => 
        \CoreAPB3_0_APBmslave0_PADDR_0[3]\, C => 
        \CoreTimer_0/N_151\, Y => \CoreTimer_0/DataOut_1_sqmuxa\);
    
    \RD_pad[6]/U0/U0\ : IOPAD_TRI
      port map(D => \RD_pad[6]/U0/NET1\, E => \RD_pad[6]/U0/NET2\, 
        PAD => RD(6));
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_24\ : NOR3C
      port map(A => \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, B => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[24]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[24]\);
    
    \CoreTimer_0/un5_intclren_0_a3_0_a2\ : NOR2
      port map(A => \CoreAPB3_0_APBmslave0_PADDR[3]\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, Y => 
        \CoreTimer_0.N_258\);
    
    \Intro_0/MSS_ADLIB_INST/U_81\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[17]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[18]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[19]INT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_41\ : MSS_IF
      port map(PIN4 => \Intro_0_MSS_MASTER_APB_PRDATA[14]\, PIN5
         => \Intro_0_MSS_MASTER_APB_PRDATA[13]\, PIN6 => 
        \Intro_0_MSS_MASTER_APB_PRDATA[15]\, PIN1 => 
        \CoreAPB3_0_APBmslave0_PWDATA[13]\, PIN2 => 
        \CoreAPB3_0_APBmslave0_PWDATA[14]\, PIN3 => 
        \CoreAPB3_0_APBmslave0_PWDATA[15]\, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[14]INT_NET\, PIN5INT
         => \Intro_0/MSS_ADLIB_INST/MSSPRDATA[13]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/MSSPRDATA[15]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[13]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[14]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[15]INT_NET\);
    
    \Intro_0/MSS_CCC_0/I_MSSCCC/U_MSSCCC\ : MSS_CCC_IP
      generic map(VCOFREQUENCY => 160.0)

      port map(CLKA => \Intro_0/MSS_CCC_0/N_CLKA_RCOSC\, EXTFB
         => \Intro_0/MSS_CCC_0/I_MSSCCC/EXTFB_INT\, GLA => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/GLA_INT\, GLAMSS => 
        \Intro_0/GLA0\, LOCK => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/LOCK_INT\, LOCKMSS => 
        \Intro_0/MSS_ADLIB_INST_PLLLOCK\, CLKB => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/CLKB_INT\, GLB => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/GLB_INT\, YB => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/YB_INT\, CLKC => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/CLKC_INT\, GLC => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/GLC_INT\, YC => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/YC_INT\, MACCLK => OPEN, SDIN
         => \Intro_0/MSS_CCC_0/I_MSSCCC/SDIN_INT\, SCLK => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/SCLK_INT\, SSHIFT => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/SSHIFT_INT\, SUPDATE => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/SUPDATE_INT\, MODE => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/MODE_INT\, SDOUT => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/SDOUT_INT\, PLLEN => 
        PLLEN_VCC, OADIV(4) => GLMUXINT_GND, OADIV(3) => 
        GLMUXINT_GND, OADIV(2) => PLLEN_VCC, OADIV(1) => 
        GLMUXINT_GND, OADIV(0) => GLMUXINT_GND, OADIVHALF => 
        GLMUXINT_GND, OADIVRST => GLMUXINT_GND, OAMUX(2) => 
        PLLEN_VCC, OAMUX(1) => GLMUXINT_GND, OAMUX(0) => 
        GLMUXINT_GND, BYPASSA => GLMUXINT_GND, DLYGLA(4) => 
        GLMUXINT_GND, DLYGLA(3) => GLMUXINT_GND, DLYGLA(2) => 
        GLMUXINT_GND, DLYGLA(1) => GLMUXINT_GND, DLYGLA(0) => 
        GLMUXINT_GND, DLYGLAMSS(4) => GLMUXINT_GND, DLYGLAMSS(3)
         => PLLEN_VCC, DLYGLAMSS(2) => GLMUXINT_GND, DLYGLAMSS(1)
         => GLMUXINT_GND, DLYGLAMSS(0) => GLMUXINT_GND, 
        DLYGLAFAB(4) => GLMUXINT_GND, DLYGLAFAB(3) => PLLEN_VCC, 
        DLYGLAFAB(2) => PLLEN_VCC, DLYGLAFAB(1) => PLLEN_VCC, 
        DLYGLAFAB(0) => PLLEN_VCC, OBDIV(4) => GLMUXINT_GND, 
        OBDIV(3) => GLMUXINT_GND, OBDIV(2) => GLMUXINT_GND, 
        OBDIV(1) => GLMUXINT_GND, OBDIV(0) => GLMUXINT_GND, 
        OBDIVHALF => GLMUXINT_GND, OBDIVRST => GLMUXINT_GND, 
        OBMUX(2) => GLMUXINT_GND, OBMUX(1) => GLMUXINT_GND, 
        OBMUX(0) => GLMUXINT_GND, BYPASSB => PLLEN_VCC, DLYGLB(4)
         => GLMUXINT_GND, DLYGLB(3) => GLMUXINT_GND, DLYGLB(2)
         => GLMUXINT_GND, DLYGLB(1) => GLMUXINT_GND, DLYGLB(0)
         => GLMUXINT_GND, OCDIV(4) => GLMUXINT_GND, OCDIV(3) => 
        GLMUXINT_GND, OCDIV(2) => GLMUXINT_GND, OCDIV(1) => 
        GLMUXINT_GND, OCDIV(0) => GLMUXINT_GND, OCDIVHALF => 
        GLMUXINT_GND, OCDIVRST => GLMUXINT_GND, OCMUX(2) => 
        GLMUXINT_GND, OCMUX(1) => GLMUXINT_GND, OCMUX(0) => 
        GLMUXINT_GND, BYPASSC => PLLEN_VCC, DLYGLC(4) => 
        GLMUXINT_GND, DLYGLC(3) => GLMUXINT_GND, DLYGLC(2) => 
        GLMUXINT_GND, DLYGLC(1) => GLMUXINT_GND, DLYGLC(0) => 
        GLMUXINT_GND, FINDIV(6) => GLMUXINT_GND, FINDIV(5) => 
        GLMUXINT_GND, FINDIV(4) => PLLEN_VCC, FINDIV(3) => 
        GLMUXINT_GND, FINDIV(2) => GLMUXINT_GND, FINDIV(1) => 
        PLLEN_VCC, FINDIV(0) => PLLEN_VCC, FBDIV(6) => 
        GLMUXINT_GND, FBDIV(5) => GLMUXINT_GND, FBDIV(4) => 
        PLLEN_VCC, FBDIV(3) => PLLEN_VCC, FBDIV(2) => PLLEN_VCC, 
        FBDIV(1) => PLLEN_VCC, FBDIV(0) => PLLEN_VCC, FBDLY(4)
         => GLMUXINT_GND, FBDLY(3) => GLMUXINT_GND, FBDLY(2) => 
        GLMUXINT_GND, FBDLY(1) => GLMUXINT_GND, FBDLY(0) => 
        PLLEN_VCC, FBSEL(1) => GLMUXINT_GND, FBSEL(0) => 
        PLLEN_VCC, XDLYSEL => GLMUXINT_GND, VCOSEL(2) => 
        GLMUXINT_GND, VCOSEL(1) => GLMUXINT_GND, VCOSEL(0) => 
        GLMUXINT_GND, GLMUXINT => GLMUXINT_GND, GLMUXSEL(1) => 
        GLMUXINT_GND, GLMUXSEL(0) => GLMUXINT_GND, GLMUXCFG(1)
         => GLMUXINT_GND, GLMUXCFG(0) => GLMUXINT_GND);
    
    \CoreTimer_0/iPRDATA_RNO_0[21]\ : MX2
      port map(A => \CoreTimer_0/Load[21]_net_1\, B => 
        \CoreTimer_0/Count[21]_net_1\, S => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, Y => 
        \CoreTimer_0/iPRDATA_RNO_0[21]_net_1\);
    
    \CoreTimer_0/Count_RNO[9]\ : AX1B
      port map(A => \CoreTimer_0/Count_c8\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_192\, Y
         => \CoreTimer_0/Count_RNO[9]_net_1\);
    
    \CoreTimer_0/PreScale_RNO[0]\ : NOR2
      port map(A => \CoreTimer_0/N_16_2\, B => 
        \CoreTimer_0/PreScale[0]_net_1\, Y => \CoreTimer_0/N_141\);
    
    \CoreTimer_0/PreScale[7]\ : DFN1C0
      port map(D => \CoreTimer_0/N_18\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => \CoreTimer_0/PreScale[7]_net_1\);
    
    \CoreTimer_0/Count_RNO[13]\ : AX1B
      port map(A => \CoreTimer_0/Count_c12\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_200\, Y
         => \CoreTimer_0/Count_RNO[13]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_94\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/I2C0SMBALERTNIINT_NET\, PIN5INT
         => \Intro_0/MSS_ADLIB_INST/I2C0BCLKINT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/I2C0SMBUSNIINT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/SPI1SSO[4]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/SPI1SSO[5]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/I2C0SMBALERTNOINT_NET\);
    
    \CoreTimer_0/PreScale_RNIT4U1[2]\ : OR2
      port map(A => \CoreTimer_0/PreScale_i_0[2]\, B => 
        \CoreTimer_0/N_144\, Y => \CoreTimer_0/N_145\);
    
    \CoreTimer_0/iPRDATA[31]\ : DFN1C0
      port map(D => \CoreTimer_0/PrdataNext[31]\, CLK => FAB_CLK, 
        CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[31]\);
    
    \CoreTimer_0/iPRDATA[0]\ : DFN1C0
      port map(D => \CoreTimer_0/N_25\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[0]\);
    
    \CoreTimer_0/iPRDATA_RNO_3[2]\ : NOR3A
      port map(A => \CoreAPB3_0_APBmslave0_PADDR_0[2]\, B => 
        \CoreAPB3_0_APBmslave0_PADDR_0[3]\, C => 
        \CoreTimer_0/Count[2]_net_1\, Y => \CoreTimer_0/N_237\);
    
    \CoreTimer_0/CtrlReg[2]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[2]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un6_ctrlen_0_a2_0_a2_net_1\, Q => 
        \CoreTimer_0/CtrlReg[2]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO_3[1]\ : NOR3A
      port map(A => \CoreAPB3_0_APBmslave0_PADDR_0[2]\, B => 
        \CoreAPB3_0_APBmslave0_PADDR_0[3]\, C => 
        \CoreTimer_0/Count[1]_net_1\, Y => 
        \CoreTimer_0/iPRDATA_RNO_3[1]_net_1\);
    
    \CoreTimer_0/Count_RNO_0[27]\ : MX2
      port map(A => \CoreTimer_0/Count[27]_net_1\, B => 
        \CoreTimer_0/Load[27]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_228\);
    
    \CoreTimer_0/iPRDATA[3]\ : DFN1C0
      port map(D => \CoreTimer_0/N_131\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[3]\);
    
    \RD_pad[0]/U0/U0\ : IOPAD_TRI
      port map(D => \RD_pad[0]/U0/NET1\, E => \RD_pad[0]/U0/NET2\, 
        PAD => RD(0));
    
    \CoreTimer_0/PreScale_RNO_0[4]\ : AO1
      port map(A => \CoreTimer_0/PreScale_i_0[4]\, B => 
        \CoreTimer_0/N_146\, C => \CoreTimer_0/LoadEnReg_net_1\, 
        Y => \CoreTimer_0/PreScale_n4_i_0_0\);
    
    \CoreTimer_0/iPRDATA_RNO[11]\ : AO1
      port map(A => \CoreTimer_0/DataOut_1_sqmuxa\, B => 
        \CoreTimer_0/Count[11]_net_1\, C => 
        \CoreTimer_0/Load_m[11]\, Y => 
        \CoreTimer_0/PrdataNext[11]\);
    
    \CoreTimer_0/Count_RNO[14]\ : AX1B
      port map(A => \CoreTimer_0/un1_loadenreg\, B => 
        \CoreTimer_0/Count_c13\, C => \CoreTimer_0/N_202\, Y => 
        \CoreTimer_0/N_381\);
    
    \FlashLED_control_wrapper_0/M1/Write_REGs.un5_wen_3\ : NOR3
      port map(A => \CoreAPB3_0_APBmslave0_PADDR[7]\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[6]\, C => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, Y => 
        \FlashLED_control_wrapper_0/M1/un5_wen_3\);
    
    \Intro_0/MSS_SPI_0_DO\ : IOPAD_TRI
      port map(D => \Intro_0/MSS_SPI_0_DO_D\, E => 
        \Intro_0/MSS_SPI_0_DO_E\, PAD => SPI_0_DO);
    
    \Intro_0/MSS_ADLIB_INST/U_72\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => \Intro_0/MSS_ADLIB_INST/FABSDD1DINT_NET\, 
        PIN5INT => \Intro_0/MSS_ADLIB_INST/FABSDD0DINT_NET\, 
        PIN6INT => OPEN, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/CMP3INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/CMP4INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/CMP5INT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_7\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/UART0CTSnINT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/GPI[31]INT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/UART0DSRnINT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/GPO[31]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/SPI0SSO[1]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/SPI0SSO[2]INT_NET\);
    
    \FlashLED_control_wrapper_0/M1/REG_control_RNIJQVQ3[0]\ : 
        NOR3B
      port map(A => \FlashLED_control_wrapper_0/M1/un2_rwclk_5\, 
        B => \FlashLED_control_wrapper_0/M1/un2_rwclk_4\, C => 
        FAB_CLK, Y => \FlashLED_control_wrapper_0/M1/un2_rwclk\);
    
    \FlashLED_control_wrapper_0/M1/RD[0]\ : DLN1
      port map(D => 
        \FlashLED_control_wrapper_0/M1/REG_load_value[0]_net_1\, 
        G => \FlashLED_control_wrapper_0/M1/un2_rwclk\, Q => 
        \RD_c[0]\);
    
    \CoreTimer_0/TimerPre_RNIILUR[1]\ : NOR2
      port map(A => \CoreTimer_0/TimerPre[1]_net_1\, B => 
        \CoreTimer_0/TimerPre[3]_net_1\, Y => 
        \CoreTimer_0/N_480_1\);
    
    \CoreTimer_0/iPRDATA_RNO[31]\ : AO1
      port map(A => \CoreTimer_0/DataOut_1_sqmuxa\, B => 
        \CoreTimer_0/Count[31]_net_1\, C => 
        \CoreTimer_0/Load_m[31]\, Y => 
        \CoreTimer_0/PrdataNext[31]\);
    
    \CoreTimer_0/CountPulse_RNO_2\ : NOR2A
      port map(A => \CoreTimer_0/PreScale[9]_net_1\, B => 
        \CoreTimer_0/N_441\, Y => \CoreTimer_0/N_482\);
    
    \CoreTimer_0/Count_RNI1RBK5[17]\ : OR2
      port map(A => \CoreTimer_0/Count_c16\, B => 
        \CoreTimer_0/Count[17]_net_1\, Y => 
        \CoreTimer_0/Count_c17\);
    
    \CoreTimer_0/iPRDATA_RNO_0[3]\ : NOR2A
      port map(A => \CoreAPB3_0_APBmslave0_PADDR[3]\, B => 
        \CoreTimer_0/TimerPre[3]_net_1\, Y => \CoreTimer_0/N_245\);
    
    \CoreTimer_0/Count_RNIC5S61[23]\ : OR3
      port map(A => \CoreTimer_0/Count[23]_net_1\, B => 
        \CoreTimer_0/Count[9]_net_1\, C => 
        \CoreTimer_0/N_58_i_0_o2_8\, Y => 
        \CoreTimer_0/N_58_i_0_o2_18\);
    
    \CoreTimer_0/CountPulse_RNO_8\ : NOR3B
      port map(A => \CoreTimer_0/PreScale[0]_net_1\, B => 
        \CoreTimer_0/N_480_1\, C => 
        \CoreTimer_0/TimerPre[2]_net_1\, Y => 
        \CoreTimer_0/NextCountPulse_0_0_a3_2_1\);
    
    \CoreTimer_0/iPRDATA_RNO_6[0]\ : NOR2A
      port map(A => \CoreAPB3_0_APBmslave0_PADDR[4]\, B => 
        \CoreTimer_0/RawTimInt_net_1\, Y => \CoreTimer_0/N_487\);
    
    \CoreTimer_0/iPRDATA_RNO_0[22]\ : MX2
      port map(A => \CoreTimer_0/Load[22]_net_1\, B => 
        \CoreTimer_0/Count[22]_net_1\, S => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, Y => 
        \CoreTimer_0/iPRDATA_RNO_0[22]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_93\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/I2C0SMBUSNOINT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/I2C1SMBUSNOINT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/CALIBOUTINT_NET\);
    
    \CoreTimer_0/Load[22]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[22]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\, Q => 
        \CoreTimer_0/Load[22]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO_2[0]\ : OR3
      port map(A => \CoreTimer_0/N_487\, B => \CoreTimer_0/N_492\, 
        C => \CoreTimer_0/N_485\, Y => 
        \CoreTimer_0/PrdataNext_iv_0_i_4[0]\);
    
    \Intro_0/MSS_ADLIB_INST/U_77\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[5]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[6]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[7]INT_NET\);
    
    \CoreTimer_0/Count[20]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[20]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte_0\, Q => 
        \CoreTimer_0/Count[20]_net_1\);
    
    \CoreTimer_0/Count[11]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[11]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte_0\, Q => 
        \CoreTimer_0/Count[11]_net_1\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_3\ : NOR3C
      port map(A => \CoreAPB3_0.iPSELS_raw_0[1]\, B => 
        \CoreAPB3_0.iPSELS_raw_1[1]\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[3]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[3]\);
    
    \CoreTimer_0/Load[21]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[21]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\, Q => 
        \CoreTimer_0/Load[21]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO_10[0]\ : OR2B
      port map(A => \CoreTimer_0/CtrlReg[1]_net_1\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, Y => 
        \CoreTimer_0/N_448\);
    
    \Intro_0/MSS_ADLIB_INST/U_91\ : MSS_IF
      port map(PIN4 => FAB_CLK, PIN5 => GLMUXINT_GND, PIN6 => 
        GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => OPEN, 
        PIN4INT => \Intro_0/MSS_ADLIB_INST/SYNCCLKFDBKINT_NET\, 
        PIN5INT => OPEN, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[31]INT_NET\, PIN1INT
         => \Intro_0/MSS_ADLIB_INST/FABPRDATA[31]INT_NET\, 
        PIN2INT => GLMUXINT_GND, PIN3INT => GLMUXINT_GND);
    
    \CoreTimer_0/iPRDATA[17]\ : DFN1C0
      port map(D => \CoreTimer_0/PrdataNext[17]\, CLK => FAB_CLK, 
        CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[17]\);
    
    \CoreTimer_0/Count_RNO_0[11]\ : MX2
      port map(A => \CoreTimer_0/Count[11]_net_1\, B => 
        \CoreTimer_0/Load[11]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_196\);
    
    \FlashLED_control_wrapper_0/M1/REG_control[3]\ : DLN1
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[3]\, G => 
        \FlashLED_control_wrapper_0/M1/REG_control_0_sqmuxa_net_1\, 
        Q => \FlashLED_control_wrapper_0/M1/REG_control[3]_net_1\);
    
    \CoreTimer_0/Load[10]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[10]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0\, Q => 
        \CoreTimer_0/Load[10]_net_1\);
    
    \CoreTimer_0/iPRDATA[25]\ : DFN1C0
      port map(D => \CoreTimer_0/PrdataNext[25]\, CLK => FAB_CLK, 
        CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[25]\);
    
    \CoreTimer_0/PreScale_RNITC91[1]\ : OR2B
      port map(A => \CoreTimer_0/PreScale[1]_net_1\, B => 
        \CoreTimer_0/PreScale[0]_net_1\, Y => \CoreTimer_0/N_144\);
    
    \Intro_0/MSS_ADLIB_INST_RNIK7F/U_CLKSRC\ : CLKSRC
      port map(A => \Intro_0/MSS_ADLIB_INST_M2FRESETn\, Y => 
        Intro_0_M2F_RESET_N);
    
    \FlashLED_control_wrapper_0/M1/RD[1]\ : DLN1
      port map(D => 
        \FlashLED_control_wrapper_0/M1/REG_load_value[1]_net_1\, 
        G => \FlashLED_control_wrapper_0/M1/un2_rwclk\, Q => 
        \RD_c[1]\);
    
    \CoreTimer_0/Count_RNO_0[9]\ : MX2
      port map(A => \CoreTimer_0/Count[9]_net_1\, B => 
        \CoreTimer_0/Load[9]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_192\);
    
    \Intro_0/MSS_ADLIB_INST/U_64\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => \Intro_0/MSS_ADLIB_INST/LVTTL4ENINT_NET\, 
        PIN5INT => \Intro_0/MSS_ADLIB_INST/LVTTL3ENINT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/LVTTL5ENINT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/LVTTL3INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/LVTTL4INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/LVTTL5INT_NET\);
    
    \CoreTimer_0/iPRDATA_RNO_2[1]\ : AO1A
      port map(A => \CoreTimer_0/CtrlReg[1]_net_1\, B => 
        \CoreTimer_0/N_257\, C => 
        \CoreTimer_0/iPRDATA_RNO_3[1]_net_1\, Y => 
        \CoreTimer_0/PrdataNext_0_iv_0_i_1[1]\);
    
    \CoreTimer_0/Count_RNO_0[15]\ : MX2
      port map(A => \CoreTimer_0/Count[15]_net_1\, B => 
        \CoreTimer_0/Load[15]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_204\);
    
    \CoreTimer_0/PreScale[4]\ : DFN1P0
      port map(D => \CoreTimer_0/N_24\, CLK => FAB_CLK, PRE => 
        Intro_0_M2F_RESET_N, Q => \CoreTimer_0/PreScale_i_0[4]\);
    
    \CoreTimer_0/iPRDATA[4]\ : DFN1C0
      port map(D => \CoreTimer_0/PrdataNext[4]\, CLK => FAB_CLK, 
        CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[4]\);
    
    \FlashLED_control_wrapper_0/M1/Write_REGs.un5_wen_1\ : NOR2
      port map(A => \CoreAPB3_0_APBmslave0_PADDR[0]\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, Y => 
        \FlashLED_control_wrapper_0/M1/un5_wen_1\);
    
    \CoreTimer_0/iPRDATA[26]\ : DFN1C0
      port map(D => \CoreTimer_0/PrdataNext[26]\, CLK => FAB_CLK, 
        CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[26]\);
    
    \CoreTimer_0/Count_RNO_1[31]\ : MX2
      port map(A => \CoreTimer_0/Count[31]_net_1\, B => 
        \CoreTimer_0/Load[31]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_236\);
    
    \CoreTimer_0/iPRDATA_RNO_0[23]\ : NOR2B
      port map(A => \CoreTimer_0/DataOut_0_sqmuxa\, B => 
        \CoreTimer_0/Load[23]_net_1\, Y => 
        \CoreTimer_0/Load_m[23]\);
    
    \Intro_0/MSS_ADLIB_INST_RNIK7F_1\ : BUFF
      port map(A => \CoreAPB3_0_APBmslave0_PADDR[3]\, Y => 
        \CoreAPB3_0_APBmslave0_PADDR_0[3]\);
    
    \FlashLED_control_wrapper_0/M1/REG_control_RNI9STS[2]\ : NOR2
      port map(A => 
        \FlashLED_control_wrapper_0/M1/REG_control[2]_net_1\, B
         => \FlashLED_control_wrapper_0/M1/REG_control[3]_net_1\, 
        Y => \FlashLED_control_wrapper_0/M1/un2_rwclk_1\);
    
    \CoreTimer_0/Count_RNO_0[20]\ : MX2
      port map(A => \CoreTimer_0/Count[20]_net_1\, B => 
        \CoreTimer_0/Load[20]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_214\);
    
    \RD_pad[1]/U0/U0\ : IOPAD_TRI
      port map(D => \RD_pad[1]/U0/NET1\, E => \RD_pad[1]/U0/NET2\, 
        PAD => RD(1));
    
    \CoreTimer_0/Count_RNIIG7D7[23]\ : OR2
      port map(A => \CoreTimer_0/Count[23]_net_1\, B => 
        \CoreTimer_0/Count_c22\, Y => \CoreTimer_0/Count_c23\);
    
    \CoreTimer_0/CountPulse_RNO_4\ : OA1C
      port map(A => \CoreTimer_0/TimerPre[0]_net_1\, B => 
        \CoreTimer_0/PreScale[7]_net_1\, C => 
        \CoreTimer_0/TimerPre[3]_net_1\, Y => 
        \CoreTimer_0/NextCountPulse_0_0_a3_0\);
    
    \CoreTimer_0/iPRDATA[29]\ : DFN1C0
      port map(D => \CoreTimer_0/N_123\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[29]\);
    
    \CoreTimer_0/TimerPre[1]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[1]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_prescaleen_0_a2_1_a3_net_1\, Q => 
        \CoreTimer_0/TimerPre[1]_net_1\);
    
    \CoreTimer_0/Count_RNO[6]\ : AX1B
      port map(A => \CoreTimer_0/Count_c5\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_186\, Y
         => \CoreTimer_0/Count_RNO[6]_net_1\);
    
    \CoreTimer_0/Count_RNITIPE2[13]\ : OR3
      port map(A => \CoreTimer_0/N_58_i_0_o2_6\, B => 
        \CoreTimer_0/N_58_i_0_o2_5\, C => 
        \CoreTimer_0/N_58_i_0_o2_18\, Y => 
        \CoreTimer_0/N_58_i_0_o2_23\);
    
    \CoreTimer_0/CountPulse_RNO_12\ : NOR2
      port map(A => \CoreTimer_0/TimerPre[3]_net_1\, B => 
        \CoreTimer_0/TimerPre[2]_net_1\, Y => 
        \CoreTimer_0/NextCountPulse_0_0_a3_0_0\);
    
    \FlashLED_control_wrapper_0/M1/Write_REGs.un5_wen\ : NOR3C
      port map(A => \FlashLED_control_wrapper_0/M1/un5_wen_2\, B
         => \FlashLED_control_wrapper_0/M1/un5_wen_1\, C => 
        \FlashLED_control_wrapper_0/M1/un5_wen_3\, Y => 
        \FlashLED_control_wrapper_0/M1/un5_wen\);
    
    \RD_pad[5]/U0/U0\ : IOPAD_TRI
      port map(D => \RD_pad[5]/U0/NET1\, E => \RD_pad[5]/U0/NET2\, 
        PAD => RD(5));
    
    \Intro_0/MSS_ADLIB_INST/U_32\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => 
        \CoreAPB3_0_APBmslave0_PADDR[6]\, PIN2 => 
        \CoreAPB3_0_APBmslave0_PADDR[7]\, PIN3 => 
        \Intro_0_MSS_MASTER_APB_PADDR[8]\, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[7]INT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[6]INT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[8]INT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[6]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[7]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[8]INT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_3\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => \Intro_0/MSS_ADLIB_INST/GPI[20]INT_NET\, 
        PIN5INT => \Intro_0/MSS_ADLIB_INST/GPI[19]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/GPI[21]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/GPO[19]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/GPO[20]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/GPO[21]INT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_10\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => \Intro_0/MSS_ADLIB_INST/VRONINT_NET\, 
        PIN5INT => \Intro_0/MSS_ADLIB_INST/RXEVINT_NET\, PIN6INT
         => \Intro_0/MSS_ADLIB_INST/CALIBININT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/UART1RTSnINT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/UART1DTRnINT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/TXEVINT_NET\);
    
    \CoreTimer_0/iPRDATA_RNO[27]\ : AO1
      port map(A => \CoreTimer_0/DataOut_1_sqmuxa\, B => 
        \CoreTimer_0/Count[27]_net_1\, C => 
        \CoreTimer_0/Load_m[27]\, Y => 
        \CoreTimer_0/PrdataNext[27]\);
    
    \Intro_0/MSS_ADLIB_INST/U_63\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/VCC15GOODINT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/VCC33GOODINT_NET\, 
        PIN3INT => GLMUXINT_GND);
    
    \CoreTimer_0/Count_RNO_1[0]\ : NOR2B
      port map(A => \CoreTimer_0/un1_loadenreg\, B => 
        \CoreTimer_0/Counte\, Y => 
        \CoreTimer_0/Count_RNO_1[0]_net_1\);
    
    \CoreTimer_0/Load[24]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[24]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\, Q => 
        \CoreTimer_0/Load[24]_net_1\);
    
    \CoreTimer_0/Count[24]\ : DFN1E1P0
      port map(D => \CoreTimer_0/N_391\, CLK => FAB_CLK, PRE => 
        Intro_0_M2F_RESET_N, E => \CoreTimer_0/Counte_0\, Q => 
        \CoreTimer_0/Count[24]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO[0]\ : NOR3
      port map(A => \CoreTimer_0/N_486\, B => 
        \CoreTimer_0/PrdataNext_iv_0_i_3[0]\, C => 
        \CoreTimer_0/PrdataNext_iv_0_i_4[0]\, Y => 
        \CoreTimer_0/N_25\);
    
    \RD_pad[2]/U0/U0\ : IOPAD_TRI
      port map(D => \RD_pad[2]/U0/NET1\, E => \RD_pad[2]/U0/NET2\, 
        PAD => RD(2));
    
    \CoreTimer_0/IntClr_RNO_0\ : NOR2B
      port map(A => \CoreTimer_0.N_258\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, Y => 
        \CoreTimer_0/un5_intclren_0_a3_0_a3_1\);
    
    \CoreTimer_0/Count_RNO_0[23]\ : MX2
      port map(A => \CoreTimer_0/Count[23]_net_1\, B => 
        \CoreTimer_0/Load[23]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_220\);
    
    \FlashLED_control_wrapper_0/M1/REG_control[0]\ : DLN1
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[0]\, G => 
        \FlashLED_control_wrapper_0/M1/REG_control_0_sqmuxa_net_1\, 
        Q => \FlashLED_control_wrapper_0/M1/REG_control[0]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_61\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => PLLEN_VCC, PIN6 => 
        GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => OPEN, 
        PIN4INT => \Intro_0/MSS_ADLIB_INST/DMAREADY[0]INT_NET\, 
        PIN5INT => \Intro_0/MSS_ADLIB_INST/F2MRESETnINT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/DMAREADY[1]INT_NET\, 
        PIN1INT => GLMUXINT_GND, PIN2INT => GLMUXINT_GND, PIN3INT
         => GLMUXINT_GND);
    
    \CoreTimer_0/Load[26]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[26]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\, Q => 
        \CoreTimer_0/Load[26]_net_1\);
    
    \RD_pad[3]/U0/U0\ : IOPAD_TRI
      port map(D => \RD_pad[3]/U0/NET1\, E => \RD_pad[3]/U0/NET2\, 
        PAD => RD(3));
    
    \CoreTimer_0/Count_RNO[15]\ : AX1B
      port map(A => \CoreTimer_0/un1_loadenreg\, B => 
        \CoreTimer_0/Count_c14\, C => \CoreTimer_0/N_204\, Y => 
        \CoreTimer_0/N_382\);
    
    \RD_pad[4]/U0/U1\ : IOTRI_OB_EB
      port map(D => \RD_c[4]\, E => PLLEN_VCC, DOUT => 
        \RD_pad[4]/U0/NET1\, EOUT => \RD_pad[4]/U0/NET2\);
    
    \Intro_0/MSS_ADLIB_INST/U_37\ : MSS_IF
      port map(PIN4 => \Intro_0_MSS_MASTER_APB_PRDATA[2]\, PIN5
         => \Intro_0_MSS_MASTER_APB_PRDATA[1]\, PIN6 => 
        \Intro_0_MSS_MASTER_APB_PRDATA[3]\, PIN1 => 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, PIN2 => 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, PIN3 => 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[2]INT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[1]INT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[3]INT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[1]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[2]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[3]INT_NET\);
    
    \CoreTimer_0/iPRDATA_RNO_0[16]\ : MX2
      port map(A => \CoreTimer_0/Load[16]_net_1\, B => 
        \CoreTimer_0/Count[16]_net_1\, S => 
        \CoreAPB3_0_APBmslave0_PADDR_0[2]\, Y => 
        \CoreTimer_0/iPRDATA_RNO_0[16]_net_1\);
    
    \CoreTimer_0/PreScale_RNI7FH4[6]\ : OR2
      port map(A => \CoreTimer_0/PreScale_i_0[6]\, B => 
        \CoreTimer_0/N_150\, Y => \CoreTimer_0/N_152\);
    
    \CoreTimer_0/iPRDATA_RNO_1[1]\ : NOR3B
      port map(A => \CoreAPB3_0_APBmslave0_PADDR_0[3]\, B => 
        \CoreAPB3_0_APBmslave0_PADDR_0[2]\, C => 
        \CoreTimer_0/TimerPre[1]_net_1\, Y => 
        \CoreTimer_0/iPRDATA_RNO_1[1]_net_1\);
    
    \CoreTimer_0/LoadEnReg_RNI439GA\ : OR2
      port map(A => \CoreTimer_0/LoadEnReg_net_1\, B => 
        \CoreTimer_0/CtrlReg_RNIC1I6A[2]_net_1\, Y => 
        \CoreTimer_0/N_16_2\);
    
    \CoreTimer_0/iPRDATA_RNO[13]\ : AO1
      port map(A => \CoreTimer_0/DataOut_1_sqmuxa\, B => 
        \CoreTimer_0/Count[13]_net_1\, C => 
        \CoreTimer_0/Load_m[13]\, Y => 
        \CoreTimer_0/PrdataNext[13]\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_16\ : NOR3C
      port map(A => \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, B => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[16]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[16]\);
    
    \CoreTimer_0/iPRDATA_RNO_0[15]\ : NOR2B
      port map(A => \CoreTimer_0/DataOut_0_sqmuxa\, B => 
        \CoreTimer_0/Load[15]_net_1\, Y => 
        \CoreTimer_0/Load_m[15]\);
    
    \CoreTimer_0/iPRDATA_RNO[29]\ : NOR3A
      port map(A => \CoreTimer_0/N_461\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, C => 
        \CoreTimer_0/N_151\, Y => \CoreTimer_0/N_123\);
    
    \CoreTimer_0/iPRDATA[30]\ : DFN1C0
      port map(D => \CoreTimer_0/N_125\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[30]\);
    
    \CoreTimer_0/Count_RNO_0[18]\ : MX2
      port map(A => \CoreTimer_0/Count[18]_net_1\, B => 
        \CoreTimer_0/Load[18]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_210\);
    
    \Intro_0/MSS_ADLIB_INST/U_78\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[8]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[9]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[10]INT_NET\);
    
    \CoreTimer_0/iPRDATA_RNO_0[28]\ : MX2
      port map(A => \CoreTimer_0/Load[28]_net_1\, B => 
        \CoreTimer_0/Count[28]_net_1\, S => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, Y => 
        \CoreTimer_0/N_460\);
    
    \CoreTimer_0/iPRDATA_RNO[1]\ : NOR3
      port map(A => \CoreTimer_0/PrdataNext_0_iv_0_i_0[1]\, B => 
        \CoreTimer_0/iPRDATA_RNO_1[1]_net_1\, C => 
        \CoreTimer_0/PrdataNext_0_iv_0_i_1[1]\, Y => 
        \CoreTimer_0/N_29\);
    
    \Intro_0/MSS_CCC_0/I_MSSCCC/U_TILE1\ : MSS_CCC_GL_IF
      port map(PIN2 => GLMUXINT_GND, PIN3 => GLMUXINT_GND, PIN4
         => GLMUXINT_GND, PIN1 => OPEN, PIN5 => FAB_CLK, PIN2INT
         => \Intro_0/MSS_CCC_0/I_MSSCCC/EXTFB_INT\, PIN3INT => 
        OPEN, PIN4INT => OPEN, PIN1INT => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/LOCK_INT\, PIN5INT => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/GLA_INT\);
    
    \FlashLED_control_wrapper_0/M1/RD[2]\ : DLN1
      port map(D => 
        \FlashLED_control_wrapper_0/M1/REG_load_value[2]_net_1\, 
        G => \FlashLED_control_wrapper_0/M1/un2_rwclk\, Q => 
        \RD_c[2]\);
    
    \CoreTimer_0/RawTimInt\ : DFN1C0
      port map(D => \CoreTimer_0/RawTimInt_RNO_net_1\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreTimer_0/RawTimInt_net_1\);
    
    \CoreTimer_0/Count_RNIU8TI[15]\ : OR2
      port map(A => \CoreTimer_0/Count[17]_net_1\, B => 
        \CoreTimer_0/Count[15]_net_1\, Y => 
        \CoreTimer_0/N_58_i_0_o2_8\);
    
    \CoreTimer_0/iPRDATA_RNO[16]\ : NOR3A
      port map(A => \CoreTimer_0/iPRDATA_RNO_0[16]_net_1\, B => 
        \CoreAPB3_0_APBmslave0_PADDR_0[3]\, C => 
        \CoreTimer_0/N_151\, Y => \CoreTimer_0/N_105\);
    
    \CoreTimer_0/Count_RNIVDQU1[5]\ : OR2
      port map(A => \CoreTimer_0/Count_c4\, B => 
        \CoreTimer_0/Count[5]_net_1\, Y => \CoreTimer_0/Count_c5\);
    
    \CoreTimer_0/Count_RNI5TN37[22]\ : OR2
      port map(A => \CoreTimer_0/Count_c21\, B => 
        \CoreTimer_0/Count[22]_net_1\, Y => 
        \CoreTimer_0/Count_c22\);
    
    \CoreTimer_0/Count_RNI2HE15[15]\ : OR2
      port map(A => \CoreTimer_0/Count[15]_net_1\, B => 
        \CoreTimer_0/Count_c14\, Y => \CoreTimer_0/Count_c15\);
    
    \FlashLED_control_wrapper_0/M1/REG_control[1]\ : DLN1
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[1]\, G => 
        \FlashLED_control_wrapper_0/M1/REG_control_0_sqmuxa_net_1\, 
        Q => \FlashLED_control_wrapper_0/M1/REG_control[1]_net_1\);
    
    \CoreTimer_0/PreScale_RNO_0[3]\ : AO1A
      port map(A => \CoreTimer_0/PreScale[3]_net_1\, B => 
        \CoreTimer_0/N_145\, C => \CoreTimer_0/LoadEnReg_net_1\, 
        Y => \CoreTimer_0/PreScale_n3_i_0_0\);
    
    \CoreTimer_0/iPRDATA[24]\ : DFN1C0
      port map(D => \CoreTimer_0/PrdataNext[24]\, CLK => FAB_CLK, 
        CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[24]\);
    
    \CoreTimer_0/Count_RNIG86J8[27]\ : OR2
      port map(A => \CoreTimer_0/Count_c26\, B => 
        \CoreTimer_0/Count[27]_net_1\, Y => 
        \CoreTimer_0/Count_c27\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_26\ : NOR3C
      port map(A => \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, B => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[26]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[26]\);
    
    \CoreTimer_0/iPRDATA_RNO_3[0]\ : OR2A
      port map(A => \CoreTimer_0/TimerPre[0]_net_1\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, Y => 
        \CoreTimer_0/N_447\);
    
    \FlashLED_control_wrapper_0/M1/RD[3]\ : DLN1
      port map(D => 
        \FlashLED_control_wrapper_0/M1/REG_load_value[3]_net_1\, 
        G => \FlashLED_control_wrapper_0/M1/un2_rwclk\, Q => 
        \RD_c[3]\);
    
    \CoreTimer_0/Count_RNI7BHE4[13]\ : OR2
      port map(A => \CoreTimer_0/Count[13]_net_1\, B => 
        \CoreTimer_0/Count_c12\, Y => \CoreTimer_0/Count_c13\);
    
    \CoreTimer_0/PreScale_RNO[6]\ : OR3A
      port map(A => \CoreTimer_0/N_152\, B => 
        \CoreTimer_0/PreScale_n6_i_0_0\, C => 
        \CoreTimer_0/CtrlReg_RNIC1I6A[2]_net_1\, Y => 
        \CoreTimer_0/N_20\);
    
    \CoreTimer_0/Count_RNIV5KQ4[18]\ : OR3
      port map(A => \CoreTimer_0/N_58_i_0_o2_20\, B => 
        \CoreTimer_0/N_58_i_0_o2_19\, C => 
        \CoreTimer_0/N_58_i_0_o2_25\, Y => 
        \CoreTimer_0/N_58_i_0_o2_27\);
    
    \CoreTimer_0/Load[8]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[8]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0\, Q => 
        \CoreTimer_0/Load[8]_net_1\);
    
    \CoreAPB3_0/iPSELS_raw_1_0[1]\ : NOR2A
      port map(A => \Intro_0_MSS_MASTER_APB_PADDR[8]\, B => 
        \Intro_0_MSS_MASTER_APB_PADDR[9]\, Y => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\);
    
    \CoreTimer_0/un5_loaden_0_a2_2_a3\ : NOR2B
      port map(A => \CoreTimer_0/N_261\, B => \CoreTimer_0.N_258\, 
        Y => \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_30\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => 
        \CoreAPB3_0_APBmslave0_PADDR[0]\, PIN2 => 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, PIN3 => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[1]INT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[0]INT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[2]INT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[0]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[1]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[2]INT_NET\);
    
    \CoreTimer_0/PreScale_RNO_0[6]\ : AO1
      port map(A => \CoreTimer_0/PreScale_i_0[6]\, B => 
        \CoreTimer_0/N_150\, C => \CoreTimer_0/LoadEnReg_net_1\, 
        Y => \CoreTimer_0/PreScale_n6_i_0_0\);
    
    \CoreTimer_0/iPRDATA[21]\ : DFN1C0
      port map(D => \CoreTimer_0/N_117\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[21]\);
    
    \CoreTimer_0/Count_RNI9TFS[31]\ : OR3
      port map(A => \CoreTimer_0/Count[24]_net_1\, B => 
        \CoreTimer_0/Count[31]_net_1\, C => 
        \CoreTimer_0/Count[25]_net_1\, Y => 
        \CoreTimer_0/N_58_i_0_o2_14\);
    
    \Intro_0/MSS_ADLIB_INST/U_75\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => GLMUXINT_GND, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[0]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/ACEFLAGS[1]INT_NET\);
    
    \CoreTimer_0/Count_RNO_0[16]\ : MX2
      port map(A => \CoreTimer_0/Count[16]_net_1\, B => 
        \CoreTimer_0/Load[16]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_206\);
    
    \CoreTimer_0/PreScale_RNO[2]\ : OR3A
      port map(A => \CoreTimer_0/N_145\, B => 
        \CoreTimer_0/PreScale_n2_i_0_0\, C => 
        \CoreTimer_0/CtrlReg_RNIC1I6A[2]_net_1\, Y => 
        \CoreTimer_0/N_28\);
    
    \CoreTimer_0/iPRDATA_RNO_0[1]\ : AO1A
      port map(A => \CoreTimer_0/Load[1]_net_1\, B => 
        \CoreTimer_0.N_258\, C => \CoreTimer_0/N_151\, Y => 
        \CoreTimer_0/PrdataNext_0_iv_0_i_0[1]\);
    
    \CoreTimer_0/CountPulse_RNIRNFE\ : NOR2B
      port map(A => \CoreTimer_0/CountPulse_net_1\, B => 
        \CoreTimer_0/CtrlReg[0]_net_1\, Y => 
        \CoreTimer_0/Countlde_0_0_a3_0\);
    
    \CoreTimer_0/un3_prdatanexten_0_a2_0\ : NOR3B
      port map(A => \CoreAPB3_0.iPSELS_raw_0[1]\, B => 
        \CoreAPB3_0.iPSELS_raw_1[1]\, C => 
        CoreAPB3_0_APBmslave0_PENABLE, Y => \CoreTimer_0/N_102\);
    
    \CoreTimer_0/Load[9]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[9]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0\, Q => 
        \CoreTimer_0/Load[9]_net_1\);
    
    \CoreTimer_0/Load[17]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[17]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\, Q => 
        \CoreTimer_0/Load[17]_net_1\);
    
    \CoreTimer_0/PrdataNext_0_iv_0_i_o3[1]\ : OR3A
      port map(A => \CoreTimer_0/N_102\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, C => 
        CoreAPB3_0_APBmslave0_PWRITE, Y => \CoreTimer_0/N_151\);
    
    \CoreTimer_0/iPRDATA[8]\ : DFN1C0
      port map(D => \CoreTimer_0/N_37\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[8]\);
    
    \CoreTimer_0/Count_RNO_0[19]\ : MX2
      port map(A => \CoreTimer_0/Count[19]_net_1\, B => 
        \CoreTimer_0/Load[19]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_212\);
    
    \CoreTimer_0/Count_RNILQ569[29]\ : OR2
      port map(A => \CoreTimer_0/Count_c28\, B => 
        \CoreTimer_0/Count[29]_net_1\, Y => 
        \CoreTimer_0/Count_c29\);
    
    \CoreTimer_0/iPRDATA_RNO_0[10]\ : NOR2B
      port map(A => \CoreTimer_0/DataOut_0_sqmuxa\, B => 
        \CoreTimer_0/Load[10]_net_1\, Y => 
        \CoreTimer_0/Load_m[10]\);
    
    \CoreTimer_0/iPRDATA_RNO[3]\ : NOR3
      port map(A => \CoreTimer_0/N_245\, B => \CoreTimer_0/N_246\, 
        C => \CoreTimer_0/PrdataNext_0_iv_0_i_1[3]\, Y => 
        \CoreTimer_0/N_131\);
    
    \CoreTimer_0/RawTimInt_RNO_0\ : NOR2A
      port map(A => \CoreTimer_0/CountIsZeroReg_i_0\, B => 
        \CoreTimer_0/N_180\, Y => \CoreTimer_0/N_255\);
    
    \FlashLED_control_wrapper_0/M1/REG_control_1_sqmuxa\ : NOR3B
      port map(A => FAB_CLK, B => 
        \FlashLED_control_wrapper_0/M1/un2_wen_3\, C => 
        \FlashLED_control_wrapper_0/M1/un5_wen\, Y => 
        \FlashLED_control_wrapper_0/M1/REG_control_1_sqmuxa_net_1\);
    
    \CoreTimer_0/Count_RNO_0[21]\ : MX2
      port map(A => \CoreTimer_0/Count[21]_net_1\, B => 
        \CoreTimer_0/Load[21]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_216\);
    
    \CoreTimer_0/Count_RNO[3]\ : MX2A
      port map(A => \CoreTimer_0/N_191_i\, B => 
        \CoreTimer_0/Load[3]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => 
        \CoreTimer_0/Count_RNO[3]_net_1\);
    
    \CoreTimer_0/Count_RNO[0]\ : MX2
      port map(A => \CoreTimer_0/Counte_mux\, B => 
        \CoreTimer_0/Load[0]_net_1\, S => 
        \CoreTimer_0/Count_RNO_1[0]_net_1\, Y => 
        \CoreTimer_0/N_507_mux\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0\ : NOR3C
      port map(A => \CoreAPB3_0.iPSELS_raw_0[1]\, B => 
        \CoreAPB3_0.iPSELS_raw_1[1]\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[0]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[0]\);
    
    \CoreTimer_0/iPRDATA[22]\ : DFN1C0
      port map(D => \CoreTimer_0/N_119\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[22]\);
    
    \CoreTimer_0/Count[22]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[22]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte_0\, Q => 
        \CoreTimer_0/Count[22]_net_1\);
    
    \CoreTimer_0/PreScale_RNO_0[2]\ : AO1
      port map(A => \CoreTimer_0/PreScale_i_0[2]\, B => 
        \CoreTimer_0/N_144\, C => \CoreTimer_0/LoadEnReg_net_1\, 
        Y => \CoreTimer_0/PreScale_n2_i_0_0\);
    
    \CoreTimer_0/PreScale_RNI3JS3[5]\ : OR2A
      port map(A => \CoreTimer_0/PreScale[5]_net_1\, B => 
        \CoreTimer_0/N_148\, Y => \CoreTimer_0/N_150\);
    
    \RD_pad[7]/U0/U0\ : IOPAD_TRI
      port map(D => \RD_pad[7]/U0/NET1\, E => \RD_pad[7]/U0/NET2\, 
        PAD => RD(7));
    
    \CoreTimer_0/iPRDATA_RNO_0[27]\ : NOR2B
      port map(A => \CoreTimer_0/DataOut_0_sqmuxa\, B => 
        \CoreTimer_0/Load[27]_net_1\, Y => 
        \CoreTimer_0/Load_m[27]\);
    
    \CoreTimer_0/IntClr\ : DFN1P0
      port map(D => \CoreTimer_0/IntClr_RNO_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, Q => 
        \CoreTimer_0/IntClr_i_0\);
    
    \CoreTimer_0/Count_RNO[23]\ : AX1B
      port map(A => \CoreTimer_0/Count_c22\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_220\, Y
         => \CoreTimer_0/Count_RNO[23]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_56\ : MSS_IF
      port map(PIN4 => \Intro_0_MSS_MASTER_APB_PRDATA[26]\, PIN5
         => \Intro_0_MSS_MASTER_APB_PRDATA[25]\, PIN6 => 
        \Intro_0_MSS_MASTER_APB_PRDATA[27]\, PIN1 => 
        \CoreAPB3_0_APBmslave0_PWDATA[25]\, PIN2 => 
        \CoreAPB3_0_APBmslave0_PWDATA[26]\, PIN3 => 
        \CoreAPB3_0_APBmslave0_PWDATA[27]\, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[26]INT_NET\, PIN5INT
         => \Intro_0/MSS_ADLIB_INST/MSSPRDATA[25]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/MSSPRDATA[27]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[25]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[26]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[27]INT_NET\);
    
    \FlashLED_control_wrapper_0/M1/Write_REGs.un2_wen_0\ : NOR3
      port map(A => \Intro_0_MSS_MASTER_APB_PADDR[11]\, B => 
        \Intro_0_MSS_MASTER_APB_PADDR[10]\, C => 
        \Intro_0_MSS_MASTER_APB_PADDR[8]\, Y => 
        \FlashLED_control_wrapper_0/M1/un2_wen_0\);
    
    \CoreTimer_0/Load[28]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[28]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\, Q => 
        \CoreTimer_0/Load[28]_net_1\);
    
    \CoreTimer_0/Load[13]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[13]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0\, Q => 
        \CoreTimer_0/Load[13]_net_1\);
    
    \CoreTimer_0/Count_RNO_0[25]\ : MX2
      port map(A => \CoreTimer_0/Count[25]_net_1\, B => 
        \CoreTimer_0/Load[25]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_224\);
    
    \CoreTimer_0/CountPulse_RNO_7\ : AO1
      port map(A => \CoreTimer_0/NextCountPulse_0_0_a3_2_1\, B
         => \CoreTimer_0/N_440\, C => \CoreTimer_0/N_479\, Y => 
        \CoreTimer_0/NextCountPulse_0_0_0\);
    
    \CoreTimer_0/Count_RNO[12]\ : AX1B
      port map(A => \CoreTimer_0/un1_loadenreg\, B => 
        \CoreTimer_0/Count_c11\, C => \CoreTimer_0/N_198\, Y => 
        \CoreTimer_0/N_379\);
    
    \CoreTimer_0/CountPulse_RNO_1\ : AO1A
      port map(A => \CoreTimer_0/N_152\, B => 
        \CoreTimer_0/NextCountPulse_0_0_a3_0\, C => 
        \CoreTimer_0/NextCountPulse_0_0_1\, Y => 
        \CoreTimer_0/NextCountPulse_0_0_2\);
    
    \CoreTimer_0/LoadEnReg_RNI42U2A_0/U_CLKSRC\ : CLKSRC
      port map(A => \CoreTimer_0/LoadEnReg_RNI42U2A_net_1\, Y => 
        \CoreTimer_0/un1_loadenreg\);
    
    \CoreTimer_0/iPRDATA[15]\ : DFN1C0
      port map(D => \CoreTimer_0/PrdataNext[15]\, CLK => FAB_CLK, 
        CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[15]\);
    
    \CoreTimer_0/iPRDATA_RNO_2[3]\ : OR3
      port map(A => \CoreTimer_0/N_151\, B => \CoreTimer_0/N_257\, 
        C => \CoreTimer_0/N_244\, Y => 
        \CoreTimer_0/PrdataNext_0_iv_0_i_1[3]\);
    
    \CoreTimer_0/Count_RNIQ9UK[3]\ : OR2
      port map(A => \CoreTimer_0/Count[7]_net_1\, B => 
        \CoreTimer_0/Count[3]_net_1\, Y => 
        \CoreTimer_0/N_58_i_0_o2_5\);
    
    \CoreTimer_0/iPRDATA[28]\ : DFN1C0
      port map(D => \CoreTimer_0/N_121\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[28]\);
    
    \CoreTimer_0/Count_RNO[24]\ : AX1B
      port map(A => \CoreTimer_0/un1_loadenreg\, B => 
        \CoreTimer_0/Count_c23\, C => \CoreTimer_0/N_222\, Y => 
        \CoreTimer_0/N_391\);
    
    \Intro_0/MSS_ADLIB_INST/U_38\ : MSS_IF
      port map(PIN4 => \Intro_0_MSS_MASTER_APB_PRDATA[5]\, PIN5
         => \Intro_0_MSS_MASTER_APB_PRDATA[4]\, PIN6 => 
        \Intro_0_MSS_MASTER_APB_PRDATA[6]\, PIN1 => 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, PIN2 => 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, PIN3 => 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[5]INT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[4]INT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[6]INT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[4]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[5]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[6]INT_NET\);
    
    \CoreTimer_0/LoadEnReg\ : DFN1C0
      port map(D => \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\, CLK
         => FAB_CLK, CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreTimer_0/LoadEnReg_net_1\);
    
    \CoreTimer_0/Count_RNO[4]\ : AX1B
      port map(A => \CoreTimer_0/Count_c3\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_182\, Y
         => \CoreTimer_0/Count_RNO[4]_net_1\);
    
    \FlashLED_control_wrapper_0/M1/REG_load_value[2]\ : DLN1
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[2]\, G => 
        \FlashLED_control_wrapper_0/M1/REG_control_1_sqmuxa_net_1\, 
        Q => 
        \FlashLED_control_wrapper_0/M1/REG_load_value[2]_net_1\);
    
    \CoreTimer_0/Count_RNO_0[30]\ : MX2
      port map(A => \CoreTimer_0/Count[30]_net_1\, B => 
        \CoreTimer_0/Load[30]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_234\);
    
    \CoreTimer_0/un5_prescaleen_0_a2_1_a3\ : NOR3C
      port map(A => \CoreAPB3_0_APBmslave0_PADDR_0[3]\, B => 
        \CoreAPB3_0_APBmslave0_PADDR_0[2]\, C => 
        \CoreTimer_0/N_261\, Y => 
        \CoreTimer_0/un5_prescaleen_0_a2_1_a3_net_1\);
    
    \CoreTimer_0/PreScale[1]\ : DFN1C0
      port map(D => \CoreTimer_0/N_30\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => \CoreTimer_0/PreScale[1]_net_1\);
    
    \CoreTimer_0/Count_RNIC07P9[12]\ : OR3
      port map(A => \CoreTimer_0/N_58_i_0_o2_23\, B => 
        \CoreTimer_0/N_58_i_0_o2_22\, C => 
        \CoreTimer_0/N_58_i_0_o2_27\, Y => \CoreTimer_0/N_180\);
    
    \CoreTimer_0/iPRDATA[16]\ : DFN1C0
      port map(D => \CoreTimer_0/N_105\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[16]\);
    
    \CoreTimer_0/Count_RNO_0[8]\ : MX2
      port map(A => \CoreTimer_0/Count[8]_net_1\, B => 
        \CoreTimer_0/Load[8]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_190\);
    
    \CoreTimer_0/PreScale_RNO[1]\ : XA1B
      port map(A => \CoreTimer_0/PreScale[0]_net_1\, B => 
        \CoreTimer_0/PreScale[1]_net_1\, C => 
        \CoreTimer_0/N_16_2\, Y => \CoreTimer_0/N_30\);
    
    \CoreTimer_0/iPRDATA[23]\ : DFN1C0
      port map(D => \CoreTimer_0/PrdataNext[23]\, CLK => FAB_CLK, 
        CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[23]\);
    
    \CoreTimer_0/Count_RNO_0[0]\ : XOR2
      port map(A => \CoreTimer_0/Counte\, B => 
        \CoreTimer_0/Count[0]_net_1\, Y => 
        \CoreTimer_0/Counte_mux\);
    
    \CoreTimer_0/Count[15]\ : DFN1E1P0
      port map(D => \CoreTimer_0/N_382\, CLK => FAB_CLK, PRE => 
        Intro_0_M2F_RESET_N, E => \CoreTimer_0/Counte_0\, Q => 
        \CoreTimer_0/Count[15]_net_1\);
    
    \FlashLED_control_wrapper_0/M1/REG_load_value[6]\ : DLN1
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[6]\, G => 
        \FlashLED_control_wrapper_0/M1/REG_control_1_sqmuxa_net_1\, 
        Q => 
        \FlashLED_control_wrapper_0/M1/REG_load_value[6]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO_0[0]\ : NOR3C
      port map(A => \CoreAPB3_0_APBmslave0_PADDR_0[3]\, B => 
        \CoreAPB3_0_APBmslave0_PADDR_0[2]\, C => 
        \CoreTimer_0/N_447\, Y => \CoreTimer_0/N_486\);
    
    \CoreTimer_0/LoadEnReg_RNI42U2A\ : OR2A
      port map(A => \CoreTimer_0/N_180\, B => 
        \CoreTimer_0/LoadEnReg_net_1\, Y => 
        \CoreTimer_0/LoadEnReg_RNI42U2A_net_1\);
    
    \CoreTimer_0/Count_RNO[18]\ : AX1B
      port map(A => \CoreTimer_0/un1_loadenreg\, B => 
        \CoreTimer_0/Count_c17\, C => \CoreTimer_0/N_210\, Y => 
        \CoreTimer_0/N_385\);
    
    \CoreTimer_0/iPRDATA_RNO[14]\ : NOR3A
      port map(A => \CoreTimer_0/N_453\, B => 
        \CoreAPB3_0_APBmslave0_PADDR_0[3]\, C => 
        \CoreTimer_0/N_151\, Y => \CoreTimer_0/N_100\);
    
    \CoreTimer_0/Count_RNO_0[14]\ : MX2
      port map(A => \CoreTimer_0/Count[14]_net_1\, B => 
        \CoreTimer_0/Load[14]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_202\);
    
    \CoreTimer_0/Count_RNO[2]\ : AX1B
      port map(A => \CoreTimer_0/N_153\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_178\, Y
         => \CoreTimer_0/Count_RNO[2]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_79\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[11]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[12]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[13]INT_NET\);
    
    \CoreTimer_0/Count_RNO[10]\ : AX1B
      port map(A => \CoreTimer_0/Count_c9\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_194\, Y
         => \CoreTimer_0/Count_RNO[10]_net_1\);
    
    \CoreTimer_0/Count[18]\ : DFN1E1P0
      port map(D => \CoreTimer_0/N_385\, CLK => FAB_CLK, PRE => 
        Intro_0_M2F_RESET_N, E => \CoreTimer_0/Counte_0\, Q => 
        \CoreTimer_0/Count[18]_net_1\);
    
    \CoreTimer_0/iPRDATA[19]\ : DFN1C0
      port map(D => \CoreTimer_0/N_113\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[19]\);
    
    \Intro_0/MSS_ADLIB_INST/U_35\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[16]INT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[15]INT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[17]INT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[15]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[16]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[17]INT_NET\);
    
    \CoreTimer_0/PreScale_RNO[3]\ : NOR3A
      port map(A => \CoreTimer_0/N_146\, B => 
        \CoreTimer_0/PreScale_n3_i_0_0\, C => 
        \CoreTimer_0/CtrlReg_RNIC1I6A[2]_net_1\, Y => 
        \CoreTimer_0/N_26\);
    
    \CoreTimer_0/Count[5]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[5]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte\, Q => \CoreTimer_0/Count[5]_net_1\);
    
    \CoreTimer_0/Count[31]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[31]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte\, Q => \CoreTimer_0/Count[31]_net_1\);
    
    \CoreTimer_0/PreScale_RNO[9]\ : XA1C
      port map(A => \CoreTimer_0/N_441\, B => 
        \CoreTimer_0/PreScale[9]_net_1\, C => 
        \CoreTimer_0/N_16_2\, Y => \CoreTimer_0/N_136\);
    
    \CoreTimer_0/iPRDATA_RNO_4[0]\ : NOR3A
      port map(A => \CoreAPB3_0_APBmslave0_PADDR[2]\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, C => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, Y => 
        \CoreTimer_0/PrdataNext_iv_0_i_a3_3_0[0]\);
    
    \Intro_0/MSS_CCC_0/I_MSSCCC/U_TILE3\ : MSS_CCC_GL_IF
      port map(PIN2 => GLMUXINT_GND, PIN3 => GLMUXINT_GND, PIN4
         => GLMUXINT_GND, PIN1 => OPEN, PIN5 => OPEN, PIN2INT => 
        OPEN, PIN3INT => \Intro_0/MSS_CCC_0/I_MSSCCC/CLKC_INT\, 
        PIN4INT => \Intro_0/MSS_CCC_0/I_MSSCCC/SUPDATE_INT\, 
        PIN1INT => \Intro_0/MSS_CCC_0/I_MSSCCC/YC_INT\, PIN5INT
         => \Intro_0/MSS_CCC_0/I_MSSCCC/GLC_INT\);
    
    \CoreTimer_0/PreScale_n8_i_0_a3_0_0\ : NOR2A
      port map(A => \CoreTimer_0/un6_ctrlen_0_a2_0_a2_net_1\, B
         => \CoreAPB3_0_APBmslave0_PWDATA[2]\, Y => 
        \CoreTimer_0/PreScale_n8_i_0_a3_0_0_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO[21]\ : NOR3A
      port map(A => \CoreTimer_0/iPRDATA_RNO_0[21]_net_1\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, C => 
        \CoreTimer_0/N_151\, Y => \CoreTimer_0/N_117\);
    
    \CoreTimer_0/Count_RNIS28U2[8]\ : OR2
      port map(A => \CoreTimer_0/Count_c7\, B => 
        \CoreTimer_0/Count[8]_net_1\, Y => \CoreTimer_0/Count_c8\);
    
    \CoreTimer_0/Count_RNO_0[4]\ : MX2
      port map(A => \CoreTimer_0/Count[4]_net_1\, B => 
        \CoreTimer_0/Load[4]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_182\);
    
    \Intro_0/MSS_ADLIB_INST/U_74\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABSDD1CLKINT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/FABSDD0CLKINT_NET\, PIN6INT => 
        OPEN, PIN1INT => GLMUXINT_GND, PIN2INT => GLMUXINT_GND, 
        PIN3INT => GLMUXINT_GND);
    
    \CoreTimer_0/Load[12]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[12]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0\, Q => 
        \CoreTimer_0/Load[12]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO[12]\ : NOR3A
      port map(A => \CoreTimer_0/N_452\, B => 
        \CoreAPB3_0_APBmslave0_PADDR_0[3]\, C => 
        \CoreTimer_0/N_151\, Y => 
        \CoreTimer_0/iPRDATA_RNO[12]_net_1\);
    
    \CoreTimer_0/Count_RNIO2TI[12]\ : OR2
      port map(A => \CoreTimer_0/Count[14]_net_1\, B => 
        \CoreTimer_0/Count[12]_net_1\, Y => 
        \CoreTimer_0/N_58_i_0_o2_2\);
    
    \CoreTimer_0/iPRDATA_RNO[5]\ : AO1
      port map(A => \CoreTimer_0/DataOut_1_sqmuxa\, B => 
        \CoreTimer_0/Count[5]_net_1\, C => 
        \CoreTimer_0/Load_m[5]\, Y => \CoreTimer_0/PrdataNext[5]\);
    
    \CoreTimer_0/Count_RNO_0[28]\ : MX2
      port map(A => \CoreTimer_0/Count[28]_net_1\, B => 
        \CoreTimer_0/Load[28]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_230\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_12\ : NOR3C
      port map(A => \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, B => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[12]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[12]\);
    
    \CoreTimer_0/Load[30]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[30]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\, Q => 
        \CoreTimer_0/Load[30]_net_1\);
    
    \CoreTimer_0/Count_RNI05NM7[24]\ : OR2
      port map(A => \CoreTimer_0/Count_c23\, B => 
        \CoreTimer_0/Count[24]_net_1\, Y => 
        \CoreTimer_0/Count_c24\);
    
    \CoreTimer_0/Load[11]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[11]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0\, Q => 
        \CoreTimer_0/Load[11]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_86\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[17]INT_NET\, PIN5INT
         => \Intro_0/MSS_ADLIB_INST/FABPWDATA[16]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/FABPWDATA[18]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[16]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[17]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[18]INT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_46\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => 
        \Intro_0/MSS_ADLIB_INST_M2FRESETn\, PIN3 => OPEN, PIN4INT
         => \Intro_0/MSS_ADLIB_INST/FABPADDR[28]INT_NET\, PIN5INT
         => \Intro_0/MSS_ADLIB_INST/FABPADDR[27]INT_NET\, PIN6INT
         => \Intro_0/MSS_ADLIB_INST/FABPADDR[29]INT_NET\, PIN1INT
         => \Intro_0/MSS_ADLIB_INST/MSSINT[5]INT_NET\, PIN2INT
         => \Intro_0/MSS_ADLIB_INST/M2FRESETnINT_NET\, PIN3INT
         => \Intro_0/MSS_ADLIB_INST/MSSINT[6]INT_NET\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_31\ : NOR3C
      port map(A => \CoreAPB3_0.iPSELS_raw_0[1]\, B => 
        \CoreAPB3_0.iPSELS_raw_1[1]\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[31]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[31]\);
    
    \CoreTimer_0/iPRDATA_RNO_1[3]\ : NOR3A
      port map(A => \CoreAPB3_0_APBmslave0_PADDR_0[2]\, B => 
        \CoreAPB3_0_APBmslave0_PADDR_0[3]\, C => 
        \CoreTimer_0/Count[3]_net_1\, Y => \CoreTimer_0/N_246\);
    
    \CoreTimer_0/iPRDATA_RNO_0[19]\ : MX2
      port map(A => \CoreTimer_0/Load[19]_net_1\, B => 
        \CoreTimer_0/Count[19]_net_1\, S => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, Y => 
        \CoreTimer_0/iPRDATA_RNO_0[19]_net_1\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_22\ : NOR3C
      port map(A => \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, B => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[22]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[22]\);
    
    \FlashLED_control_wrapper_0/M1/RD[5]\ : DLN1
      port map(D => 
        \FlashLED_control_wrapper_0/M1/REG_load_value[5]_net_1\, 
        G => \FlashLED_control_wrapper_0/M1/un2_rwclk\, Q => 
        \RD_c[5]\);
    
    \CoreTimer_0/CountPulse_RNO_6\ : OA1A
      port map(A => \CoreTimer_0/TimerPre[0]_net_1\, B => 
        \CoreTimer_0/PreScale[5]_net_1\, C => 
        \CoreTimer_0/N_480_1\, Y => 
        \CoreTimer_0/NextCountPulse_0_0_a3_1_0\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_7\ : NOR3C
      port map(A => \CoreAPB3_0.iPSELS_raw_0[1]\, B => 
        \CoreAPB3_0.iPSELS_raw_1[1]\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[7]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[7]\);
    
    \Intro_0/MSS_ADLIB_INST/U_73\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/FABACETRIGINT_NET\, PIN6INT => 
        OPEN, PIN1INT => \Intro_0/MSS_ADLIB_INST/CMP6INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/CMP7INT_NET\, PIN3INT
         => GLMUXINT_GND);
    
    \CoreTimer_0/iPRDATA_RNO[15]\ : AO1
      port map(A => \CoreTimer_0/DataOut_1_sqmuxa\, B => 
        \CoreTimer_0/Count[15]_net_1\, C => 
        \CoreTimer_0/Load_m[15]\, Y => 
        \CoreTimer_0/PrdataNext[15]\);
    
    \CoreTimer_0/iPRDATA[20]\ : DFN1C0
      port map(D => \CoreTimer_0/N_115\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[20]\);
    
    \CoreTimer_0/Load[25]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[25]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\, Q => 
        \CoreTimer_0/Load[25]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO_0[30]\ : MX2
      port map(A => \CoreTimer_0/Load[30]_net_1\, B => 
        \CoreTimer_0/Count[30]_net_1\, S => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, Y => 
        \CoreTimer_0/iPRDATA_RNO_0[30]_net_1\);
    
    \CoreTimer_0/iPRDATA[14]\ : DFN1C0
      port map(D => \CoreTimer_0/N_100\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[14]\);
    
    \CoreTimer_0/Count_RNO_0[26]\ : MX2
      port map(A => \CoreTimer_0/Count[26]_net_1\, B => 
        \CoreTimer_0/Load[26]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_226\);
    
    \CoreTimer_0/Count_RNO[30]\ : AX1B
      port map(A => \CoreTimer_0/Count_c29\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_234\, Y
         => \CoreTimer_0/Count_RNO[30]_net_1\);
    
    \FlashLED_control_wrapper_0/M1/REG_load_value[3]\ : DLN1
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[3]\, G => 
        \FlashLED_control_wrapper_0/M1/REG_control_1_sqmuxa_net_1\, 
        Q => 
        \FlashLED_control_wrapper_0/M1/REG_load_value[3]_net_1\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_5\ : NOR3C
      port map(A => \CoreAPB3_0.iPSELS_raw_0[1]\, B => 
        \CoreAPB3_0.iPSELS_raw_1[1]\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[5]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[5]\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_17\ : NOR3C
      port map(A => \CoreAPB3_0/iPSELS_raw_0_0[1]_net_1\, B => 
        \CoreAPB3_0/iPSELS_raw_1_0[1]_net_1\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[17]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[17]\);
    
    \Intro_0/MSS_UART_0_RXD\ : IOPAD_IN
      port map(PAD => UART_0_RXD, Y => \Intro_0/MSS_UART_0_RXD_Y\);
    
    \CoreTimer_0/CtrlReg_RNIB5QFA[2]\ : OA1A
      port map(A => \CoreTimer_0/CtrlReg[2]_net_1\, B => 
        \CoreTimer_0/N_180\, C => \CoreTimer_0/Countlde_0_0_a3_0\, 
        Y => \CoreTimer_0/N_248\);
    
    \RD_pad[6]/U0/U1\ : IOTRI_OB_EB
      port map(D => \RD_c[6]\, E => PLLEN_VCC, DOUT => 
        \RD_pad[6]/U0/NET1\, EOUT => \RD_pad[6]/U0/NET2\);
    
    \CoreTimer_0/PreScale_RNO_0[5]\ : AO1A
      port map(A => \CoreTimer_0/PreScale[5]_net_1\, B => 
        \CoreTimer_0/N_148\, C => \CoreTimer_0/LoadEnReg_net_1\, 
        Y => \CoreTimer_0/PreScale_n5_i_0_0\);
    
    \CoreTimer_0/Count_RNIFQ608[25]\ : OR2
      port map(A => \CoreTimer_0/Count_c24\, B => 
        \CoreTimer_0/Count[25]_net_1\, Y => 
        \CoreTimer_0/Count_c25\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_30\ : NOR3C
      port map(A => \CoreAPB3_0.iPSELS_raw_0[1]\, B => 
        \CoreAPB3_0.iPSELS_raw_1[1]\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[30]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[30]\);
    
    \Intro_0/MSS_ADLIB_INST/U_71\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/CMP0INT_NET\, PIN2INT
         => \Intro_0/MSS_ADLIB_INST/CMP1INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/CMP2INT_NET\);
    
    \CoreTimer_0/Count_RNIJTSI[10]\ : OR2
      port map(A => \CoreTimer_0/Count[10]_net_1\, B => 
        \CoreTimer_0/Count[11]_net_1\, Y => 
        \CoreTimer_0/N_58_i_0_o2_13\);
    
    \CoreTimer_0/CountPulse_RNO_10\ : NOR3B
      port map(A => \CoreTimer_0/N_443\, B => 
        \CoreTimer_0/NextCountPulse_0_0_a3_0_0\, C => 
        \CoreTimer_0/N_145\, Y => \CoreTimer_0/N_479\);
    
    \CoreTimer_0/iPRDATA[11]\ : DFN1C0
      port map(D => \CoreTimer_0/PrdataNext[11]\, CLK => FAB_CLK, 
        CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[11]\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_27\ : NOR3C
      port map(A => \CoreAPB3_0.iPSELS_raw_0[1]\, B => 
        \CoreAPB3_0.iPSELS_raw_1[1]\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[27]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[27]\);
    
    \CoreTimer_0/Load[6]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[6]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0\, Q => 
        \CoreTimer_0/Load[6]_net_1\);
    
    \CoreTimer_0/Count_RNO_0[29]\ : MX2
      port map(A => \CoreTimer_0/Count[29]_net_1\, B => 
        \CoreTimer_0/Load[29]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_232\);
    
    \CoreTimer_0/LoadEnReg_RNIF830L_0\ : OR3
      port map(A => \CoreTimer_0/N_248\, B => 
        \CoreTimer_0/LoadEnReg_net_1\, C => 
        \CoreTimer_0/CtrlReg_RNIC1I6A[2]_net_1\, Y => 
        \CoreTimer_0/Counte\);
    
    \CoreTimer_0/Count[21]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[21]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte_0\, Q => 
        \CoreTimer_0/Count[21]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_39\ : MSS_IF
      port map(PIN4 => \Intro_0_MSS_MASTER_APB_PRDATA[8]\, PIN5
         => \Intro_0_MSS_MASTER_APB_PRDATA[7]\, PIN6 => 
        \Intro_0_MSS_MASTER_APB_PRDATA[9]\, PIN1 => 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, PIN2 => 
        \CoreAPB3_0_APBmslave0_PWDATA[8]\, PIN3 => 
        \CoreAPB3_0_APBmslave0_PWDATA[9]\, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[8]INT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[7]INT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[9]INT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[7]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[8]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPWDATA[9]INT_NET\);
    
    \CoreTimer_0/iPRDATA_RNO[4]\ : AO1
      port map(A => \CoreTimer_0/DataOut_1_sqmuxa\, B => 
        \CoreTimer_0/Count[4]_net_1\, C => 
        \CoreTimer_0/Load_m[4]\, Y => \CoreTimer_0/PrdataNext[4]\);
    
    \CoreTimer_0/Count[13]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[13]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte_0\, Q => 
        \CoreTimer_0/Count[13]_net_1\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_9\ : NOR3C
      port map(A => \CoreAPB3_0.iPSELS_raw_0[1]\, B => 
        \CoreAPB3_0.iPSELS_raw_1[1]\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[9]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[9]\);
    
    \CoreTimer_0/Count_RNO_0[31]\ : OR2
      port map(A => \CoreTimer_0/Count[30]_net_1\, B => 
        \CoreTimer_0/un1_loadenreg\, Y => 
        \CoreTimer_0/Count_66_0\);
    
    \CoreTimer_0/Count_RNO[25]\ : AX1B
      port map(A => \CoreTimer_0/un1_loadenreg\, B => 
        \CoreTimer_0/Count_c24\, C => \CoreTimer_0/N_224\, Y => 
        \CoreTimer_0/N_392\);
    
    \CoreTimer_0/Count[19]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[19]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte_0\, Q => 
        \CoreTimer_0/Count[19]_net_1\);
    
    \RD_pad[0]/U0/U1\ : IOTRI_OB_EB
      port map(D => \RD_c[0]\, E => PLLEN_VCC, DOUT => 
        \RD_pad[0]/U0/NET1\, EOUT => \RD_pad[0]/U0/NET2\);
    
    \CoreTimer_0/PreScale_RNO[8]\ : OR3A
      port map(A => \CoreTimer_0/N_441\, B => \CoreTimer_0/N_463\, 
        C => \CoreTimer_0/N_16_2\, Y => \CoreTimer_0/N_16\);
    
    \CoreTimer_0/iPRDATA_RNO_0[14]\ : MX2
      port map(A => \CoreTimer_0/Load[14]_net_1\, B => 
        \CoreTimer_0/Count[14]_net_1\, S => 
        \CoreAPB3_0_APBmslave0_PADDR_0[2]\, Y => 
        \CoreTimer_0/N_453\);
    
    \CoreTimer_0/Count_RNO_0[12]\ : MX2
      port map(A => \CoreTimer_0/Count[12]_net_1\, B => 
        \CoreTimer_0/Load[12]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_198\);
    
    \Intro_0/MSS_CCC_0/I_MSSCCC/U_TILE0\ : MSS_CCC_IF
      port map(PIN2 => GLMUXINT_GND, PIN3 => GLMUXINT_GND, PIN4
         => GLMUXINT_GND, PIN1 => OPEN, PIN2INT => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/SDIN_INT\, PIN3INT => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/SCLK_INT\, PIN4INT => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/SSHIFT_INT\, PIN1INT => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/SDOUT_INT\);
    
    \FlashLED_control_wrapper_0/M1/REG_control_0_sqmuxa\ : NOR3C
      port map(A => FAB_CLK, B => 
        \FlashLED_control_wrapper_0/M1/un2_wen_3\, C => 
        \FlashLED_control_wrapper_0/M1/un5_wen\, Y => 
        \FlashLED_control_wrapper_0/M1/REG_control_0_sqmuxa_net_1\);
    
    \CoreTimer_0/Count_RNO[8]\ : AX1B
      port map(A => \CoreTimer_0/Count_c7\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_190\, Y
         => \CoreTimer_0/Count_RNO[8]_net_1\);
    
    \CoreTimer_0/Count[9]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[9]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte\, Q => \CoreTimer_0/Count[9]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_52\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[14]INT_NET\, PIN5INT
         => \Intro_0/MSS_ADLIB_INST/FABPWDATA[13]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/FABPWDATA[15]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[13]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[14]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/FABPRDATA[15]INT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_5\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => \Intro_0/MSS_ADLIB_INST/GPI[26]INT_NET\, 
        PIN5INT => \Intro_0/MSS_ADLIB_INST/GPI[25]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/GPI[27]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/GPO[25]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/GPO[26]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/GPO[27]INT_NET\);
    
    \CoreTimer_0/Load[14]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[14]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0\, Q => 
        \CoreTimer_0/Load[14]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_34\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[13]INT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[12]INT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[14]INT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[12]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[13]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[14]INT_NET\);
    
    \CoreTimer_0/un5_prescaleen_0_a2_1_a2\ : NOR3B
      port map(A => \CoreTimer_0/N_102\, B => 
        CoreAPB3_0_APBmslave0_PWRITE, C => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, Y => 
        \CoreTimer_0/N_261\);
    
    \CoreTimer_0/iPRDATA[12]\ : DFN1C0
      port map(D => \CoreTimer_0/iPRDATA_RNO[12]_net_1\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[12]\);
    
    \CoreTimer_0/Count_RNO_0[3]\ : XOR2
      port map(A => \CoreTimer_0/N_154\, B => 
        \CoreTimer_0/Count[3]_net_1\, Y => \CoreTimer_0/N_191_i\);
    
    \Intro_0/MSS_CCC_0/I_MSSCCC/U_TILE2\ : MSS_CCC_GL_IF
      port map(PIN2 => GLMUXINT_GND, PIN3 => GLMUXINT_GND, PIN4
         => GLMUXINT_GND, PIN1 => OPEN, PIN5 => OPEN, PIN2INT => 
        OPEN, PIN3INT => \Intro_0/MSS_CCC_0/I_MSSCCC/CLKB_INT\, 
        PIN4INT => \Intro_0/MSS_CCC_0/I_MSSCCC/MODE_INT\, PIN1INT
         => \Intro_0/MSS_CCC_0/I_MSSCCC/YB_INT\, PIN5INT => 
        \Intro_0/MSS_CCC_0/I_MSSCCC/GLB_INT\);
    
    \CoreTimer_0/Count_RNI1CTI[16]\ : OR2
      port map(A => \CoreTimer_0/Count[16]_net_1\, B => 
        \CoreTimer_0/Count[19]_net_1\, Y => 
        \CoreTimer_0/N_58_i_0_o2_10\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_1\ : NOR3C
      port map(A => \CoreAPB3_0.iPSELS_raw_0[1]\, B => 
        \CoreAPB3_0.iPSELS_raw_1[1]\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[1]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[1]\);
    
    \CoreTimer_0/PreScale[5]\ : DFN1C0
      port map(D => \CoreTimer_0/N_22\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => \CoreTimer_0/PreScale[5]_net_1\);
    
    \CoreTimer_0/Count_RNISQOJ2[7]\ : OR2
      port map(A => \CoreTimer_0/Count_c6\, B => 
        \CoreTimer_0/Count[7]_net_1\, Y => \CoreTimer_0/Count_c7\);
    
    \CoreTimer_0/Load[16]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[16]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0\, Q => 
        \CoreTimer_0/Load[16]_net_1\);
    
    \CoreTimer_0/Count_RNIPA8Q6[21]\ : OR2
      port map(A => \CoreTimer_0/Count_c20\, B => 
        \CoreTimer_0/Count[21]_net_1\, Y => 
        \CoreTimer_0/Count_c21\);
    
    \CoreTimer_0/Count_RNO_0[1]\ : XOR2
      port map(A => \CoreTimer_0/Count[1]_net_1\, B => 
        \CoreTimer_0/Count[0]_net_1\, Y => \CoreTimer_0/N_190_i\);
    
    \Intro_0/MSS_CCC_0/I_RCOSC\ : RCOSC
      port map(CLKOUT => \Intro_0/MSS_CCC_0/N_CLKA_RCOSC\);
    
    \CoreAPB3_0/u_mux_p_to_b3/PRDATA_2\ : NOR3C
      port map(A => \CoreAPB3_0.iPSELS_raw_0[1]\, B => 
        \CoreAPB3_0.iPSELS_raw_1[1]\, C => 
        \CoreAPB3_0_APBmslave1_PRDATA[2]\, Y => 
        \Intro_0_MSS_MASTER_APB_PRDATA[2]\);
    
    \FlashLED_control_wrapper_0/M1/REG_control[6]\ : DLN1
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[6]\, G => 
        \FlashLED_control_wrapper_0/M1/REG_control_0_sqmuxa_net_1\, 
        Q => \FlashLED_control_wrapper_0/M1/REG_control[6]_net_1\);
    
    \CoreTimer_0/Count_RNITJR51[18]\ : OR3
      port map(A => \CoreTimer_0/Count[21]_net_1\, B => 
        \CoreTimer_0/Count[18]_net_1\, C => 
        \CoreTimer_0/N_58_i_0_o2_10\, Y => 
        \CoreTimer_0/N_58_i_0_o2_19\);
    
    \Intro_0/MSS_ADLIB_INST/U_57\ : MSS_IF
      port map(PIN4 => \Intro_0_MSS_MASTER_APB_PRDATA[29]\, PIN5
         => \Intro_0_MSS_MASTER_APB_PRDATA[28]\, PIN6 => 
        \Intro_0_MSS_MASTER_APB_PRDATA[30]\, PIN1 => 
        \CoreAPB3_0_APBmslave0_PWDATA[28]\, PIN2 => 
        \CoreAPB3_0_APBmslave0_PWDATA[29]\, PIN3 => 
        \CoreAPB3_0_APBmslave0_PWDATA[30]\, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPRDATA[29]INT_NET\, PIN5INT
         => \Intro_0/MSS_ADLIB_INST/MSSPRDATA[28]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/MSSPRDATA[30]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[28]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[29]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/MSSPWDATA[30]INT_NET\);
    
    \CoreTimer_0/CountIsZeroReg\ : DFN1P0
      port map(D => \CoreTimer_0/N_180\, CLK => FAB_CLK, PRE => 
        Intro_0_M2F_RESET_N, Q => 
        \CoreTimer_0/CountIsZeroReg_i_0\);
    
    \FlashLED_control_wrapper_0/M1/REG_control[5]\ : DLN1
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[5]\, G => 
        \FlashLED_control_wrapper_0/M1/REG_control_0_sqmuxa_net_1\, 
        Q => \FlashLED_control_wrapper_0/M1/REG_control[5]_net_1\);
    
    \CoreTimer_0/Count_RNO[19]\ : AX1B
      port map(A => \CoreTimer_0/Count_c18\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_212\, Y
         => \CoreTimer_0/Count_RNO[19]_net_1\);
    
    \CoreTimer_0/Count[17]\ : DFN1E1P0
      port map(D => \CoreTimer_0/N_384\, CLK => FAB_CLK, PRE => 
        Intro_0_M2F_RESET_N, E => \CoreTimer_0/Counte_0\, Q => 
        \CoreTimer_0/Count[17]_net_1\);
    
    \CoreTimer_0/Count_RNIG7PF2[12]\ : OR3
      port map(A => \CoreTimer_0/N_58_i_0_o2_2\, B => 
        \CoreTimer_0/N_58_i_0_o2_1\, C => 
        \CoreTimer_0/N_58_i_0_o2_16\, Y => 
        \CoreTimer_0/N_58_i_0_o2_22\);
    
    \CoreTimer_0/iPRDATA[18]\ : DFN1C0
      port map(D => \CoreTimer_0/N_110\, CLK => FAB_CLK, CLR => 
        Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[18]\);
    
    \Intro_0/MSS_ADLIB_INST/U_33\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => 
        \Intro_0_MSS_MASTER_APB_PADDR[9]\, PIN2 => 
        \Intro_0_MSS_MASTER_APB_PADDR[10]\, PIN3 => 
        \Intro_0_MSS_MASTER_APB_PADDR[11]\, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[10]INT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[9]INT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[11]INT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[9]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[10]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[11]INT_NET\);
    
    \CoreTimer_0/Load[7]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[7]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0\, Q => 
        \CoreTimer_0/Load[7]_net_1\);
    
    \CoreTimer_0/Count_RNIH0UK[1]\ : OR2
      port map(A => \CoreTimer_0/Count[0]_net_1\, B => 
        \CoreTimer_0/Count[1]_net_1\, Y => \CoreTimer_0/N_153\);
    
    \CoreTimer_0/Load[5]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[5]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0\, Q => 
        \CoreTimer_0/Load[5]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO[18]\ : NOR3A
      port map(A => \CoreTimer_0/N_455\, B => 
        \CoreAPB3_0_APBmslave0_PADDR_0[3]\, C => 
        \CoreTimer_0/N_151\, Y => \CoreTimer_0/N_110\);
    
    \CoreTimer_0/Count_RNO_0[24]\ : MX2
      port map(A => \CoreTimer_0/Count[24]_net_1\, B => 
        \CoreTimer_0/Load[24]_net_1\, S => 
        \CoreTimer_0/un1_loadenreg\, Y => \CoreTimer_0/N_222\);
    
    \CoreTimer_0/Load[1]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[1]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0\, Q => 
        \CoreTimer_0/Load[1]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO[23]\ : AO1
      port map(A => \CoreTimer_0/DataOut_1_sqmuxa\, B => 
        \CoreTimer_0/Count[23]_net_1\, C => 
        \CoreTimer_0/Load_m[23]\, Y => 
        \CoreTimer_0/PrdataNext[23]\);
    
    \CoreTimer_0/Count_RNIM2VI[20]\ : OR2
      port map(A => \CoreTimer_0/Count[20]_net_1\, B => 
        \CoreTimer_0/Count[22]_net_1\, Y => 
        \CoreTimer_0/N_58_i_0_o2_12\);
    
    \FlashLED_control_wrapper_0/M1/REG_load_value[7]\ : DLN1
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[7]\, G => 
        \FlashLED_control_wrapper_0/M1/REG_control_1_sqmuxa_net_1\, 
        Q => 
        \FlashLED_control_wrapper_0/M1/REG_load_value[7]_net_1\);
    
    \CoreTimer_0/Count_RNI21MS8[28]\ : OR2
      port map(A => \CoreTimer_0/Count_c27\, B => 
        \CoreTimer_0/Count[28]_net_1\, Y => 
        \CoreTimer_0/Count_c28\);
    
    \CoreTimer_0/iPRDATA[13]\ : DFN1C0
      port map(D => \CoreTimer_0/PrdataNext[13]\, CLK => FAB_CLK, 
        CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[13]\);
    
    \CoreTimer_0/Count_RNITJ992[6]\ : OR2
      port map(A => \CoreTimer_0/Count_c5\, B => 
        \CoreTimer_0/Count[6]_net_1\, Y => \CoreTimer_0/Count_c6\);
    
    \CoreTimer_0/iPRDATA_RNO[26]\ : AO1
      port map(A => \CoreTimer_0/DataOut_1_sqmuxa\, B => 
        \CoreTimer_0/Count[26]_net_1\, C => 
        \CoreTimer_0/Load_m[26]\, Y => 
        \CoreTimer_0/PrdataNext[26]\);
    
    \CoreTimer_0/iPRDATA_RNO[10]\ : AO1
      port map(A => \CoreTimer_0/DataOut_1_sqmuxa\, B => 
        \CoreTimer_0/Count[10]_net_1\, C => 
        \CoreTimer_0/Load_m[10]\, Y => 
        \CoreTimer_0/PrdataNext[10]\);
    
    \Intro_0/MSS_ADLIB_INST/U_31\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, PIN2 => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, PIN3 => 
        \CoreAPB3_0_APBmslave0_PADDR[5]\, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[4]INT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[3]INT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/FABPADDR[5]INT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[3]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[4]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPADDR[5]INT_NET\);
    
    \CoreTimer_0/iPRDATA_RNO[30]\ : NOR3A
      port map(A => \CoreTimer_0/iPRDATA_RNO_0[30]_net_1\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, C => 
        \CoreTimer_0/N_151\, Y => \CoreTimer_0/N_125\);
    
    \CoreTimer_0/Load[29]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[29]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_loaden_0_a2_2_a3_net_1\, Q => 
        \CoreTimer_0/Load[29]_net_1\);
    
    \FlashLED_control_wrapper_0/M1/REG_load_value[1]\ : DLN1
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[1]\, G => 
        \FlashLED_control_wrapper_0/M1/REG_control_1_sqmuxa_net_1\, 
        Q => 
        \FlashLED_control_wrapper_0/M1/REG_load_value[1]_net_1\);
    
    \CoreTimer_0/Count[16]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[16]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte_0\, Q => 
        \CoreTimer_0/Count[16]_net_1\);
    
    \CoreTimer_0/TimerPre[0]\ : DFN1E1C0
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[0]\, CLK => 
        FAB_CLK, CLR => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/un5_prescaleen_0_a2_1_a3_net_1\, Q => 
        \CoreTimer_0/TimerPre[0]_net_1\);
    
    \CoreTimer_0/RawTimInt_RNO\ : OA1
      port map(A => \CoreTimer_0/RawTimInt_net_1\, B => 
        \CoreTimer_0/N_255\, C => \CoreTimer_0/IntClr_i_0\, Y => 
        \CoreTimer_0/RawTimInt_RNO_net_1\);
    
    \CoreTimer_0/PreScale_RNIUTI2[3]\ : OR2A
      port map(A => \CoreTimer_0/PreScale[3]_net_1\, B => 
        \CoreTimer_0/N_145\, Y => \CoreTimer_0/N_146\);
    
    \RD_pad[1]/U0/U1\ : IOTRI_OB_EB
      port map(D => \RD_c[1]\, E => PLLEN_VCC, DOUT => 
        \RD_pad[1]/U0/NET1\, EOUT => \RD_pad[1]/U0/NET2\);
    
    \FlashLED_control_wrapper_0/M1/Write_REGs.un5_wen_2\ : NOR2A
      port map(A => \CoreTimer_0.N_258\, B => 
        \CoreAPB3_0_APBmslave0_PADDR[5]\, Y => 
        \FlashLED_control_wrapper_0/M1/un5_wen_2\);
    
    \CoreTimer_0/iPRDATA_RNO_0[11]\ : NOR2B
      port map(A => \CoreTimer_0/DataOut_0_sqmuxa\, B => 
        \CoreTimer_0/Load[11]_net_1\, Y => 
        \CoreTimer_0/Load_m[11]\);
    
    \Intro_0/MSS_ADLIB_INST/U_50\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[8]INT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[7]INT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWDATA[9]INT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[7]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[8]INT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/FABPRDATA[9]INT_NET\);
    
    \CoreTimer_0/iPRDATA_RNO_0[5]\ : NOR2B
      port map(A => \CoreTimer_0/DataOut_0_sqmuxa\, B => 
        \CoreTimer_0/Load[5]_net_1\, Y => \CoreTimer_0/Load_m[5]\);
    
    \CoreTimer_0/Count[8]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[8]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte\, Q => \CoreTimer_0/Count[8]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_66\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => \Intro_0/MSS_ADLIB_INST/LVTTL7ENINT_NET\, 
        PIN5INT => \Intro_0/MSS_ADLIB_INST/LVTTL6ENINT_NET\, 
        PIN6INT => OPEN, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/LVTTL6INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/LVTTL7INT_NET\, PIN3INT => 
        GLMUXINT_GND);
    
    \CoreTimer_0/Count[1]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[1]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte\, Q => \CoreTimer_0/Count[1]_net_1\);
    
    \RD_pad[5]/U0/U1\ : IOTRI_OB_EB
      port map(D => \RD_c[5]\, E => PLLEN_VCC, DOUT => 
        \RD_pad[5]/U0/NET1\, EOUT => \RD_pad[5]/U0/NET2\);
    
    \FlashLED_control_wrapper_0/M1/REG_control[2]\ : DLN1
      port map(D => \CoreAPB3_0_APBmslave0_PWDATA[2]\, G => 
        \FlashLED_control_wrapper_0/M1/REG_control_0_sqmuxa_net_1\, 
        Q => \FlashLED_control_wrapper_0/M1/REG_control[2]_net_1\);
    
    \CoreTimer_0/iPRDATA_RNO[7]\ : AO1
      port map(A => \CoreTimer_0/DataOut_1_sqmuxa\, B => 
        \CoreTimer_0/Count[7]_net_1\, C => 
        \CoreTimer_0/Load_m[7]\, Y => \CoreTimer_0/PrdataNext[7]\);
    
    \CoreTimer_0/Count_RNO[22]\ : AX1B
      port map(A => \CoreTimer_0/Count_c21\, B => 
        \CoreTimer_0/un1_loadenreg\, C => \CoreTimer_0/N_218\, Y
         => \CoreTimer_0/Count_RNO[22]_net_1\);
    
    \CoreTimer_0/Count[7]\ : DFN1E1P0
      port map(D => \CoreTimer_0/Count_RNO[7]_net_1\, CLK => 
        FAB_CLK, PRE => Intro_0_M2F_RESET_N, E => 
        \CoreTimer_0/Counte\, Q => \CoreTimer_0/Count[7]_net_1\);
    
    \Intro_0/MSS_ADLIB_INST/U_82\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => OPEN, PIN5INT => OPEN, PIN6INT => OPEN, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[20]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[21]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/ACEFLAGS[22]INT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_8\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/UART0DCDnINT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/UART0RInINT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/UART1CTSnINT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/SPI0SSO[3]INT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/UART0RTSnINT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/UART0DTRnINT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_42\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => Intro_0_MSS_MASTER_APB_PSELx, 
        PIN2 => CoreAPB3_0_APBmslave0_PENABLE, PIN3 => 
        CoreAPB3_0_APBmslave0_PWRITE, PIN4INT => 
        \Intro_0/MSS_ADLIB_INST/FABPENABLEINT_NET\, PIN5INT => 
        \Intro_0/MSS_ADLIB_INST/FABPSELINT_NET\, PIN6INT => 
        \Intro_0/MSS_ADLIB_INST/FABPWRITEINT_NET\, PIN1INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPSELINT_NET\, PIN2INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPENABLEINT_NET\, PIN3INT => 
        \Intro_0/MSS_ADLIB_INST/MSSPWRITEINT_NET\);
    
    \Intro_0/MSS_ADLIB_INST/U_4\ : MSS_IF
      port map(PIN4 => GLMUXINT_GND, PIN5 => GLMUXINT_GND, PIN6
         => GLMUXINT_GND, PIN1 => OPEN, PIN2 => OPEN, PIN3 => 
        OPEN, PIN4INT => \Intro_0/MSS_ADLIB_INST/GPI[23]INT_NET\, 
        PIN5INT => \Intro_0/MSS_ADLIB_INST/GPI[22]INT_NET\, 
        PIN6INT => \Intro_0/MSS_ADLIB_INST/GPI[24]INT_NET\, 
        PIN1INT => \Intro_0/MSS_ADLIB_INST/GPO[22]INT_NET\, 
        PIN2INT => \Intro_0/MSS_ADLIB_INST/GPO[23]INT_NET\, 
        PIN3INT => \Intro_0/MSS_ADLIB_INST/GPO[24]INT_NET\);
    
    \CoreTimer_0/iPRDATA[7]\ : DFN1C0
      port map(D => \CoreTimer_0/PrdataNext[7]\, CLK => FAB_CLK, 
        CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[7]\);
    
    \CoreTimer_0/iPRDATA[6]\ : DFN1C0
      port map(D => \CoreTimer_0/PrdataNext[6]\, CLK => FAB_CLK, 
        CLR => Intro_0_M2F_RESET_N, Q => 
        \CoreAPB3_0_APBmslave1_PRDATA[6]\);
    
    \CoreTimer_0/DataOut_0_sqmuxa_0_a2_0_a3\ : NOR3
      port map(A => \CoreAPB3_0_APBmslave0_PADDR[3]\, B => 
        \CoreTimer_0/N_151\, C => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, Y => 
        \CoreTimer_0/DataOut_0_sqmuxa\);
    
    \CoreTimer_0/PreScale_RNO_0[8]\ : OA1A
      port map(A => \CoreTimer_0/PreScale[7]_net_1\, B => 
        \CoreTimer_0/N_152\, C => \CoreTimer_0/PreScale_i_0[8]\, 
        Y => \CoreTimer_0/N_463\);
    
    \RD_pad[2]/U0/U1\ : IOTRI_OB_EB
      port map(D => \RD_c[2]\, E => PLLEN_VCC, DOUT => 
        \RD_pad[2]/U0/NET1\, EOUT => \RD_pad[2]/U0/NET2\);
    
    GND_power_inst1 : GND
      port map( Y => GND_power_net1);

    VCC_power_inst1 : VCC
      port map( Y => VCC_power_net1);


end DEF_ARCH; 
