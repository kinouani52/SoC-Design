----------------------------------------------------------------------
-- Created by Microsemi SmartDesign Tue Dec 08 09:10:13 2020
-- Parameters for CoreTimer
----------------------------------------------------------------------


LIBRARY ieee;
   USE ieee.std_logic_1164.all;
   USE ieee.std_logic_unsigned.all;
   USE ieee.numeric_std.all;

package coreparameters is
    constant FAMILY : integer := 18;
    constant INTACTIVEH : integer := 1;
    constant WIDTH : integer := 32;
end coreparameters;
